library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity bios_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of bios_rom is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"ED",X"77",X"F8",X"50",X"30",X"E8",X"4D",X"49",X"4E",X"45",X"80",X"F8",X"50",X"00",X"DE",X"53",
		X"54",X"4F",X"52",X"4D",X"80",X"00",X"8E",X"C8",X"83",X"6F",X"80",X"8C",X"CB",X"BB",X"26",X"F9",
		X"BD",X"E8",X"E3",X"7C",X"C8",X"24",X"86",X"BB",X"B7",X"C8",X"80",X"8E",X"01",X"01",X"BF",X"C8",
		X"81",X"8E",X"C8",X"83",X"6F",X"80",X"8C",X"CB",X"70",X"26",X"F9",X"20",X"00",X"BD",X"F1",X"AF",
		X"CC",X"02",X"00",X"BD",X"F7",X"A9",X"0A",X"79",X"0F",X"56",X"0F",X"9B",X"8E",X"C8",X"A8",X"BD",
		X"F8",X"4F",X"8E",X"C8",X"AF",X"BD",X"F8",X"4F",X"8E",X"C8",X"F9",X"BD",X"F8",X"4F",X"CC",X"00",
		X"01",X"BD",X"F8",X"7C",X"8E",X"C9",X"00",X"BD",X"F8",X"4F",X"CC",X"00",X"01",X"BD",X"F8",X"7C",
		X"8E",X"CB",X"B3",X"9F",X"C4",X"8E",X"CB",X"B7",X"9F",X"C6",X"C6",X"08",X"8E",X"CB",X"B3",X"BD",
		X"F5",X"3F",X"86",X"05",X"97",X"D9",X"97",X"DA",X"97",X"DB",X"20",X"23",X"BD",X"E8",X"66",X"10",
		X"8E",X"C8",X"C4",X"96",X"9B",X"AE",X"A6",X"BD",X"ED",X"AB",X"8E",X"ED",X"A7",X"96",X"9B",X"AE",
		X"86",X"A6",X"05",X"84",X"03",X"26",X"02",X"0C",X"D9",X"CC",X"00",X"01",X"BD",X"F8",X"7C",X"BD",
		X"E7",X"E4",X"8E",X"C8",X"C4",X"96",X"9B",X"AE",X"86",X"BD",X"E1",X"29",X"20",X"3B",X"DC",X"F0",
		X"83",X"00",X"01",X"DD",X"F0",X"27",X"26",X"34",X"08",X"BD",X"F1",X"AA",X"BD",X"EA",X"CF",X"CE",
		X"EE",X"2F",X"BD",X"EA",X"9D",X"35",X"08",X"8E",X"C8",X"A8",X"CE",X"CB",X"EB",X"BD",X"F8",X"D8",
		X"8E",X"C8",X"AF",X"CE",X"CB",X"EB",X"BD",X"F8",X"D8",X"96",X"0F",X"27",X"0C",X"DC",X"F0",X"10",
		X"26",X"FF",X"3E",X"7E",X"EF",X"CC",X"12",X"12",X"12",X"34",X"08",X"BD",X"EA",X"F0",X"BD",X"E5",
		X"1E",X"BD",X"E2",X"62",X"BD",X"E4",X"B8",X"BD",X"E3",X"53",X"35",X"08",X"BD",X"EB",X"43",X"BD",
		X"EC",X"46",X"BD",X"EC",X"95",X"BD",X"E6",X"47",X"25",X"DF",X"96",X"BD",X"10",X"27",X"FF",X"6C",
		X"96",X"BE",X"10",X"26",X"FF",X"98",X"7E",X"E0",X"AF",X"9F",X"C2",X"CC",X"7F",X"00",X"DD",X"DC",
		X"97",X"B7",X"86",X"20",X"97",X"9C",X"8E",X"E1",X"E7",X"9F",X"9D",X"8E",X"C9",X"33",X"9F",X"B9",
		X"86",X"1D",X"97",X"B8",X"0F",X"56",X"CE",X"ED",X"77",X"BD",X"F6",X"8D",X"34",X"08",X"BD",X"E7",
		X"11",X"BD",X"F6",X"87",X"96",X"26",X"85",X"01",X"26",X"02",X"0A",X"B7",X"BD",X"EA",X"F0",X"BD",
		X"EA",X"CF",X"BD",X"F2",X"89",X"BD",X"E5",X"1E",X"BD",X"F2",X"A5",X"F6",X"C8",X"B7",X"27",X"1C",
		X"8E",X"EF",X"26",X"10",X"BE",X"C8",X"DC",X"BD",X"EA",X"7F",X"8E",X"EF",X"5D",X"BD",X"EA",X"7F",
		X"8E",X"EF",X"94",X"BD",X"EA",X"7F",X"35",X"08",X"0A",X"DC",X"20",X"C0",X"35",X"08",X"0F",X"9C",
		X"86",X"04",X"97",X"B7",X"86",X"7F",X"97",X"B8",X"96",X"B7",X"27",X"4A",X"D6",X"B8",X"27",X"04",
		X"0A",X"B8",X"20",X"12",X"D6",X"26",X"C4",X"1F",X"26",X"0C",X"4A",X"97",X"B7",X"9E",X"C2",X"A6",
		X"86",X"C6",X"03",X"BD",X"E9",X"A1",X"34",X"08",X"BD",X"EA",X"F0",X"BD",X"F2",X"A9",X"CE",X"EE",
		X"20",X"BD",X"EA",X"9D",X"10",X"8E",X"E0",X"00",X"CE",X"ED",X"A7",X"B6",X"C8",X"9B",X"EE",X"C6",
		X"BD",X"EA",X"A8",X"BD",X"E5",X"1E",X"BD",X"E2",X"62",X"BD",X"E4",X"B8",X"35",X"08",X"BD",X"EB",
		X"43",X"BD",X"E6",X"47",X"20",X"B2",X"39",X"0A",X"B8",X"27",X"4E",X"0C",X"ED",X"BD",X"F5",X"17",
		X"84",X"07",X"8B",X"04",X"97",X"9C",X"DE",X"B9",X"86",X"80",X"A7",X"C4",X"DC",X"DC",X"8B",X"08",
		X"A7",X"44",X"6F",X"45",X"E7",X"46",X"6F",X"47",X"BD",X"F5",X"17",X"4D",X"2B",X"0C",X"81",X"10",
		X"2C",X"02",X"8B",X"0C",X"81",X"60",X"2F",X"0E",X"20",X"EE",X"81",X"F0",X"2F",X"02",X"80",X"0C",
		X"81",X"A0",X"2C",X"02",X"20",X"E2",X"A7",X"C8",X"11",X"1F",X"89",X"1D",X"8A",X"01",X"A7",X"C8",
		X"10",X"6F",X"42",X"31",X"C8",X"12",X"10",X"9F",X"B9",X"39",X"00",X"02",X"07",X"10",X"00",X"20",
		X"18",X"10",X"01",X"00",X"05",X"00",X"03",X"25",X"07",X"50",X"00",X"00",X"01",X"00",X"00",X"35",
		X"00",X"00",X"00",X"00",X"04",X"04",X"08",X"08",X"0D",X"0D",X"EE",X"3D",X"EE",X"53",X"EE",X"6F",
		X"EE",X"8E",X"34",X"08",X"86",X"C8",X"1F",X"8B",X"96",X"BD",X"10",X"26",X"00",X"9C",X"96",X"EE",
		X"10",X"26",X"00",X"A7",X"96",X"13",X"10",X"26",X"00",X"92",X"96",X"14",X"27",X"32",X"96",X"D4",
		X"91",X"D6",X"27",X"1C",X"91",X"D8",X"27",X"08",X"96",X"D5",X"27",X"14",X"96",X"D7",X"26",X"20",
		X"96",X"D7",X"8B",X"0C",X"81",X"7F",X"22",X"18",X"97",X"D7",X"96",X"D4",X"97",X"D8",X"20",X"0E",
		X"96",X"D5",X"8B",X"0C",X"81",X"7F",X"22",X"08",X"97",X"D5",X"96",X"D4",X"97",X"D6",X"0C",X"F2",
		X"96",X"D5",X"27",X"0E",X"80",X"02",X"97",X"D5",X"D6",X"D6",X"BD",X"E7",X"B5",X"10",X"9F",X"CC",
		X"9F",X"CE",X"96",X"D7",X"27",X"0E",X"80",X"02",X"97",X"D7",X"D6",X"D8",X"BD",X"E7",X"B5",X"10",
		X"9F",X"D0",X"9F",X"D2",X"DC",X"C8",X"D3",X"CC",X"D3",X"D0",X"DD",X"C8",X"DC",X"CA",X"D3",X"CE",
		X"D3",X"D2",X"DD",X"CA",X"96",X"1B",X"27",X"0F",X"2B",X"04",X"0A",X"D4",X"20",X"06",X"0C",X"D4",
		X"20",X"02",X"34",X"08",X"BD",X"E8",X"4C",X"86",X"D0",X"1F",X"8B",X"BD",X"F2",X"A5",X"C6",X"0C",
		X"10",X"8E",X"C8",X"C8",X"8E",X"CB",X"89",X"BD",X"EA",X"8D",X"35",X"88",X"86",X"80",X"97",X"EE",
		X"BD",X"F5",X"17",X"84",X"03",X"8B",X"03",X"97",X"EF",X"0C",X"F6",X"96",X"EE",X"2A",X"19",X"0A",
		X"EF",X"27",X"0D",X"BD",X"E9",X"8A",X"97",X"C8",X"0F",X"C9",X"D7",X"CA",X"0F",X"CB",X"35",X"88",
		X"04",X"EE",X"86",X"1F",X"97",X"EF",X"35",X"88",X"D6",X"EF",X"C1",X"E0",X"2F",X"0C",X"96",X"EF",
		X"80",X"04",X"97",X"EF",X"4F",X"BD",X"E9",X"4A",X"35",X"88",X"0F",X"EF",X"0F",X"EE",X"BD",X"E8",
		X"37",X"35",X"88",X"B6",X"C8",X"E7",X"27",X"2B",X"34",X"08",X"86",X"C8",X"1F",X"8B",X"12",X"12",
		X"12",X"12",X"DC",X"DE",X"D3",X"E2",X"DD",X"DE",X"97",X"DC",X"DC",X"E0",X"D3",X"E4",X"DD",X"E0",
		X"97",X"DD",X"35",X"08",X"BD",X"F2",X"A5",X"C6",X"08",X"10",X"BE",X"C8",X"DC",X"8E",X"EF",X"B3",
		X"BD",X"EA",X"7F",X"39",X"8E",X"E3",X"A1",X"9F",X"A3",X"BD",X"F5",X"17",X"8E",X"E4",X"48",X"84",
		X"06",X"AE",X"86",X"EC",X"81",X"DD",X"DC",X"97",X"DE",X"0F",X"DF",X"D7",X"E0",X"0F",X"E1",X"20",
		X"58",X"96",X"BF",X"26",X"19",X"BD",X"F5",X"17",X"84",X"7F",X"8B",X"30",X"97",X"A2",X"BD",X"F5",
		X"17",X"84",X"3F",X"97",X"E6",X"BD",X"F5",X"17",X"8B",X"10",X"97",X"E7",X"20",X"49",X"96",X"BD",
		X"26",X"E3",X"C6",X"1C",X"CE",X"C9",X"33",X"A6",X"C4",X"27",X"08",X"33",X"C8",X"12",X"5A",X"26",
		X"F6",X"20",X"34",X"0C",X"ED",X"0A",X"BF",X"9E",X"DE",X"AF",X"44",X"9E",X"E0",X"AF",X"46",X"86",
		X"40",X"A7",X"C4",X"96",X"C0",X"26",X"10",X"8E",X"E4",X"12",X"9F",X"9D",X"BD",X"F5",X"17",X"84",
		X"7F",X"8B",X"40",X"97",X"9C",X"0C",X"C0",X"9E",X"E8",X"A6",X"80",X"97",X"A2",X"A6",X"80",X"97",
		X"E6",X"A6",X"80",X"97",X"E7",X"9F",X"E8",X"D6",X"E6",X"BD",X"E7",X"B5",X"10",X"9F",X"E2",X"9F",
		X"E4",X"39",X"CE",X"C8",X"C4",X"96",X"9B",X"EE",X"C6",X"A6",X"C4",X"C6",X"03",X"BD",X"E9",X"A1",
		X"8E",X"E4",X"26",X"9F",X"9D",X"39",X"0A",X"C1",X"27",X"06",X"86",X"FF",X"97",X"9C",X"20",X"17",
		X"BD",X"F5",X"17",X"1F",X"89",X"C4",X"03",X"26",X"02",X"CB",X"01",X"CE",X"C8",X"C4",X"96",X"9B",
		X"EE",X"C6",X"A6",X"C4",X"BD",X"E9",X"A1",X"39",X"E4",X"50",X"E4",X"6A",X"E4",X"84",X"E4",X"9E",
		X"7F",X"00",X"28",X"20",X"30",X"40",X"28",X"30",X"28",X"00",X"10",X"30",X"10",X"40",X"18",X"20",
		X"50",X"40",X"30",X"28",X"30",X"08",X"60",X"7F",X"38",X"70",X"80",X"00",X"40",X"00",X"30",X"20",
		X"10",X"50",X"20",X"28",X"40",X"30",X"3E",X"70",X"18",X"30",X"60",X"20",X"18",X"40",X"30",X"24",
		X"50",X"7F",X"06",X"70",X"00",X"7F",X"40",X"10",X"60",X"28",X"38",X"30",X"28",X"08",X"40",X"30",
		X"28",X"7F",X"20",X"18",X"30",X"30",X"08",X"68",X"40",X"20",X"50",X"7F",X"38",X"70",X"00",X"80",
		X"40",X"30",X"60",X"38",X"18",X"30",X"30",X"20",X"18",X"20",X"38",X"40",X"28",X"10",X"60",X"20",
		X"00",X"30",X"40",X"38",X"50",X"7F",X"1C",X"70",X"86",X"04",X"CE",X"C9",X"0B",X"8E",X"C8",X"15",
		X"B7",X"C8",X"8F",X"BD",X"F2",X"A9",X"A6",X"C4",X"27",X"22",X"6A",X"49",X"27",X"19",X"EC",X"45",
		X"E3",X"41",X"ED",X"45",X"EC",X"47",X"E3",X"43",X"ED",X"47",X"31",X"45",X"BD",X"EA",X"6D",X"33",
		X"4A",X"7A",X"C8",X"8F",X"26",X"E0",X"39",X"6F",X"C4",X"7A",X"C8",X"EA",X"B6",X"C8",X"BD",X"26",
		X"EE",X"B6",X"C8",X"EE",X"26",X"E9",X"A6",X"84",X"27",X"E5",X"6F",X"84",X"7C",X"C8",X"B6",X"6C",
		X"C4",X"FC",X"C8",X"C8",X"ED",X"45",X"FC",X"C8",X"CA",X"ED",X"47",X"FC",X"C9",X"07",X"ED",X"41",
		X"FC",X"C9",X"09",X"ED",X"43",X"86",X"18",X"A7",X"49",X"7C",X"C8",X"EA",X"20",X"C1",X"86",X"1C",
		X"B7",X"C8",X"8F",X"CE",X"C9",X"33",X"A6",X"C4",X"26",X"09",X"33",X"C8",X"12",X"7A",X"C8",X"8F",
		X"26",X"F4",X"39",X"10",X"2B",X"00",X"9C",X"85",X"40",X"10",X"26",X"00",X"A4",X"85",X"20",X"10",
		X"26",X"00",X"A9",X"85",X"10",X"10",X"26",X"00",X"D4",X"85",X"01",X"10",X"26",X"00",X"D8",X"A6",
		X"41",X"81",X"04",X"27",X"56",X"85",X"01",X"27",X"31",X"B6",X"C8",X"EE",X"26",X"2C",X"B6",X"C8",
		X"BD",X"26",X"27",X"34",X"08",X"BD",X"F1",X"AF",X"96",X"C8",X"A0",X"44",X"D6",X"CA",X"E0",X"46",
		X"BD",X"F5",X"93",X"80",X"10",X"97",X"83",X"8E",X"E2",X"3E",X"E6",X"43",X"A6",X"85",X"D6",X"83",
		X"BD",X"E7",X"B5",X"10",X"AF",X"48",X"AF",X"4A",X"35",X"08",X"EC",X"44",X"E3",X"48",X"ED",X"44",
		X"EC",X"46",X"E3",X"4A",X"ED",X"46",X"BD",X"F2",X"A5",X"8E",X"E2",X"5A",X"A6",X"41",X"48",X"AE",
		X"86",X"31",X"44",X"E6",X"42",X"BD",X"EA",X"8D",X"7E",X"E5",X"2A",X"EC",X"44",X"E3",X"48",X"29",
		X"1A",X"ED",X"44",X"EC",X"46",X"E3",X"4A",X"29",X"12",X"ED",X"46",X"BD",X"F2",X"A9",X"31",X"44",
		X"8E",X"CB",X"A4",X"C6",X"04",X"BD",X"EA",X"8D",X"7E",X"E5",X"2A",X"6F",X"C4",X"7A",X"C8",X"EB",
		X"7E",X"E5",X"2A",X"A6",X"46",X"AB",X"C8",X"10",X"A7",X"46",X"A1",X"C8",X"11",X"26",X"02",X"64",
		X"C4",X"BD",X"F2",X"A5",X"31",X"44",X"BD",X"EA",X"6D",X"7E",X"E5",X"2A",X"A6",X"43",X"81",X"03",
		X"26",X"0D",X"A6",X"42",X"A1",X"C8",X"10",X"2C",X"06",X"8B",X"08",X"A7",X"42",X"20",X"1B",X"64",
		X"C4",X"A6",X"C8",X"10",X"A7",X"42",X"86",X"18",X"A7",X"C8",X"10",X"B6",X"C8",X"ED",X"26",X"0A",
		X"B6",X"C8",X"C0",X"26",X"05",X"86",X"7F",X"B7",X"C8",X"A2",X"7E",X"E5",X"96",X"6A",X"C8",X"10",
		X"26",X"02",X"64",X"C4",X"7E",X"E5",X"96",X"6F",X"C4",X"A6",X"41",X"81",X"04",X"27",X"15",X"E6",
		X"43",X"5A",X"27",X"10",X"34",X"0A",X"86",X"C8",X"1F",X"8B",X"A6",X"E4",X"BD",X"E9",X"A1",X"BD",
		X"E9",X"A1",X"35",X"0A",X"7E",X"E5",X"2A",X"34",X"08",X"BD",X"F1",X"AA",X"BD",X"F2",X"A9",X"CE",
		X"CB",X"2B",X"86",X"0E",X"B7",X"C8",X"8F",X"A6",X"C4",X"10",X"27",X"00",X"A6",X"E6",X"44",X"E1",
		X"41",X"24",X"0D",X"CB",X"03",X"E7",X"44",X"10",X"AE",X"42",X"8E",X"EE",X"BA",X"BD",X"EA",X"7F",
		X"4D",X"10",X"2A",X"00",X"83",X"7A",X"C8",X"F7",X"10",X"27",X"00",X"37",X"B6",X"C8",X"26",X"84",
		X"01",X"26",X"03",X"7C",X"C8",X"F8",X"B6",X"C8",X"F8",X"10",X"8E",X"7F",X"00",X"8E",X"EF",X"04",
		X"BD",X"E7",X"6A",X"10",X"8E",X"60",X"80",X"8E",X"EF",X"0B",X"BD",X"E7",X"6A",X"10",X"8E",X"80",
		X"50",X"8E",X"EF",X"15",X"BD",X"E7",X"6A",X"10",X"8E",X"A0",X"80",X"8E",X"EF",X"1C",X"BD",X"E7",
		X"6A",X"20",X"50",X"7A",X"C8",X"D9",X"7F",X"C8",X"EB",X"7F",X"C8",X"ED",X"B6",X"C8",X"79",X"27",
		X"2B",X"B6",X"C8",X"9B",X"44",X"8E",X"C8",X"DA",X"F6",X"C8",X"D9",X"E7",X"86",X"B6",X"C8",X"DA",
		X"26",X"05",X"B6",X"C8",X"DB",X"27",X"1A",X"B6",X"C8",X"9B",X"8B",X"02",X"84",X"02",X"B7",X"C8",
		X"9B",X"44",X"8E",X"C8",X"DA",X"E6",X"86",X"F7",X"C8",X"D9",X"27",X"EB",X"B6",X"C8",X"D9",X"26",
		X"0D",X"86",X"01",X"B7",X"C8",X"BE",X"20",X"06",X"E6",X"44",X"E1",X"41",X"25",X"05",X"6F",X"C4",
		X"7A",X"C8",X"EC",X"33",X"45",X"7A",X"C8",X"8F",X"10",X"26",X"FF",X"4B",X"BD",X"EC",X"C9",X"20",
		X"05",X"34",X"08",X"BD",X"F1",X"AA",X"BD",X"F2",X"A5",X"8E",X"80",X"38",X"BF",X"C8",X"90",X"BD",
		X"EF",X"D8",X"27",X"1E",X"12",X"12",X"12",X"7A",X"C8",X"8F",X"27",X"16",X"B6",X"C8",X"91",X"8B",
		X"06",X"B7",X"C8",X"91",X"C6",X"04",X"10",X"BE",X"C8",X"90",X"8E",X"EE",X"EB",X"BD",X"EA",X"7F",
		X"20",X"E5",X"35",X"08",X"96",X"26",X"84",X"01",X"48",X"48",X"48",X"8E",X"EE",X"AD",X"CE",X"CB",
		X"A4",X"BD",X"F6",X"1F",X"D6",X"EC",X"26",X"0F",X"96",X"BD",X"26",X"08",X"D6",X"EB",X"DA",X"ED",
		X"DA",X"E7",X"26",X"03",X"1C",X"FE",X"39",X"1A",X"01",X"39",X"34",X"32",X"8E",X"C8",X"C8",X"BD",
		X"F2",X"F2",X"A6",X"E4",X"97",X"04",X"1F",X"20",X"BD",X"F3",X"12",X"C6",X"0C",X"AE",X"61",X"BD",
		X"F4",X"0E",X"35",X"B2",X"34",X"16",X"8E",X"CB",X"2B",X"86",X"0E",X"E6",X"84",X"27",X"07",X"30",
		X"05",X"4A",X"26",X"F7",X"20",X"1D",X"A6",X"E4",X"84",X"80",X"4C",X"A7",X"84",X"2A",X"02",X"0C",
		X"BD",X"A6",X"E4",X"84",X"7F",X"A7",X"04",X"A6",X"61",X"A7",X"01",X"EC",X"62",X"ED",X"02",X"0C",
		X"EC",X"0C",X"F3",X"35",X"96",X"34",X"36",X"BD",X"F6",X"01",X"A7",X"64",X"1D",X"58",X"49",X"58",
		X"49",X"58",X"49",X"ED",X"62",X"E6",X"64",X"1D",X"58",X"49",X"58",X"49",X"58",X"49",X"ED",X"64",
		X"35",X"B6",X"34",X"36",X"8D",X"DF",X"EC",X"7C",X"58",X"49",X"ED",X"64",X"EC",X"7A",X"58",X"49",
		X"ED",X"62",X"35",X"B6",X"86",X"D0",X"1F",X"8B",X"BD",X"F2",X"72",X"86",X"C8",X"1F",X"8B",X"0F",
		X"9C",X"0F",X"9F",X"0F",X"A2",X"0F",X"A5",X"8E",X"C9",X"0B",X"6F",X"80",X"8C",X"CB",X"71",X"26",
		X"F9",X"CC",X"00",X"00",X"DD",X"DE",X"DD",X"E0",X"DD",X"E2",X"DD",X"E4",X"97",X"E7",X"97",X"BD",
		X"97",X"BE",X"97",X"EA",X"97",X"EB",X"97",X"EC",X"97",X"F8",X"C6",X"40",X"D7",X"F7",X"97",X"ED",
		X"97",X"C0",X"8E",X"08",X"00",X"9F",X"F0",X"86",X"07",X"97",X"BF",X"8E",X"E3",X"84",X"9F",X"A3",
		X"CC",X"00",X"00",X"DD",X"C8",X"DD",X"CA",X"CC",X"00",X"00",X"97",X"D4",X"DD",X"CC",X"DD",X"CE",
		X"97",X"D5",X"97",X"D6",X"DD",X"D0",X"DD",X"D2",X"97",X"D7",X"97",X"D8",X"96",X"D4",X"8E",X"EE",
		X"EB",X"CE",X"CB",X"89",X"BD",X"F6",X"1F",X"86",X"7F",X"D6",X"D4",X"BD",X"E7",X"D2",X"10",X"BF",
		X"C9",X"07",X"BF",X"C9",X"09",X"39",X"34",X"30",X"34",X"08",X"BD",X"F1",X"AA",X"BD",X"F2",X"72",
		X"35",X"08",X"86",X"A0",X"97",X"8F",X"96",X"C8",X"27",X"0A",X"2B",X"03",X"4A",X"20",X"01",X"4C",
		X"97",X"C8",X"0F",X"C9",X"96",X"CA",X"27",X"0A",X"2B",X"03",X"4A",X"20",X"01",X"4C",X"97",X"CA",
		X"0F",X"CB",X"96",X"D4",X"27",X"0C",X"81",X"1F",X"2E",X"03",X"4A",X"20",X"01",X"4C",X"84",X"3F",
		X"97",X"D4",X"BD",X"E2",X"F2",X"8E",X"CB",X"81",X"C6",X"08",X"A6",X"84",X"8B",X"03",X"A7",X"80",
		X"5A",X"26",X"F7",X"34",X"08",X"BD",X"F1",X"AA",X"BD",X"EA",X"CF",X"5F",X"86",X"20",X"BD",X"E9",
		X"0B",X"BD",X"E8",X"FD",X"35",X"08",X"96",X"C8",X"10",X"26",X"FF",X"AA",X"96",X"CA",X"10",X"26",
		X"FF",X"A4",X"96",X"D4",X"10",X"26",X"FF",X"9E",X"0A",X"8F",X"10",X"26",X"FF",X"98",X"BD",X"E7",
		X"E4",X"35",X"B0",X"8E",X"ED",X"E0",X"10",X"8E",X"CB",X"71",X"CE",X"CB",X"81",X"C6",X"08",X"86",
		X"16",X"AF",X"A1",X"30",X"08",X"A7",X"C0",X"8B",X"0F",X"5A",X"26",X"F5",X"39",X"34",X"1E",X"8E",
		X"CB",X"81",X"86",X"08",X"6C",X"80",X"4A",X"26",X"FB",X"20",X"02",X"34",X"1E",X"86",X"D0",X"1F",
		X"8B",X"86",X"09",X"34",X"02",X"6A",X"E4",X"26",X"07",X"BD",X"F3",X"54",X"35",X"02",X"35",X"9E",
		X"BD",X"F3",X"54",X"86",X"03",X"B7",X"C8",X"23",X"A6",X"E4",X"4A",X"8E",X"CB",X"81",X"E6",X"86",
		X"C4",X"7F",X"E1",X"61",X"23",X"DF",X"E0",X"62",X"2F",X"DB",X"D7",X"04",X"8E",X"CB",X"71",X"48",
		X"AE",X"86",X"BD",X"F2",X"A9",X"BD",X"F2",X"D5",X"20",X"CB",X"34",X"1E",X"86",X"D0",X"1F",X"8B",
		X"86",X"09",X"34",X"02",X"6A",X"E4",X"26",X"07",X"BD",X"F3",X"54",X"35",X"02",X"35",X"9E",X"BD",
		X"F3",X"54",X"86",X"03",X"B7",X"C8",X"23",X"8E",X"C8",X"C8",X"BD",X"F2",X"F2",X"E6",X"E4",X"58",
		X"58",X"EB",X"62",X"2F",X"DF",X"C4",X"7F",X"D7",X"04",X"8E",X"CB",X"71",X"A6",X"E4",X"4A",X"48",
		X"AE",X"86",X"BD",X"F2",X"A9",X"BD",X"F2",X"D5",X"20",X"CA",X"34",X"06",X"BD",X"F5",X"17",X"A7",
		X"E4",X"BD",X"F5",X"17",X"81",X"60",X"2E",X"F9",X"81",X"A0",X"2D",X"F5",X"A7",X"61",X"35",X"06",
		X"39",X"34",X"76",X"96",X"ED",X"10",X"27",X"00",X"93",X"0A",X"ED",X"BD",X"F5",X"17",X"84",X"1F",
		X"97",X"8B",X"81",X"1B",X"23",X"04",X"80",X"04",X"20",X"F6",X"C6",X"12",X"3D",X"C3",X"C9",X"33",
		X"1F",X"03",X"A6",X"C4",X"84",X"C0",X"26",X"0D",X"0C",X"8B",X"96",X"8B",X"81",X"1B",X"2F",X"EA",
		X"0F",X"8B",X"4F",X"20",X"E5",X"A6",X"E4",X"A7",X"41",X"8E",X"E2",X"42",X"48",X"10",X"AE",X"86",
		X"10",X"9F",X"89",X"C6",X"20",X"E7",X"C4",X"8E",X"E2",X"3E",X"A6",X"61",X"E6",X"86",X"D7",X"8B",
		X"8E",X"E2",X"3A",X"E6",X"86",X"E7",X"C8",X"10",X"A7",X"43",X"8E",X"E2",X"52",X"48",X"10",X"AE",
		X"86",X"10",X"AF",X"4C",X"8E",X"E2",X"4A",X"10",X"AE",X"86",X"10",X"9F",X"87",X"81",X"06",X"26",
		X"02",X"0C",X"F4",X"96",X"88",X"9B",X"8A",X"19",X"A7",X"4F",X"96",X"87",X"99",X"89",X"19",X"A7",
		X"4E",X"96",X"8B",X"BD",X"EA",X"3E",X"BD",X"E7",X"B5",X"10",X"AF",X"48",X"AF",X"4A",X"0C",X"EB",
		X"96",X"C0",X"27",X"08",X"86",X"FF",X"97",X"9C",X"86",X"03",X"97",X"C1",X"35",X"F6",X"34",X"06",
		X"BD",X"F5",X"17",X"1F",X"89",X"84",X"30",X"A7",X"61",X"C4",X"0F",X"C1",X"04",X"24",X"02",X"CB",
		X"04",X"C1",X"0C",X"23",X"02",X"C0",X"04",X"EB",X"61",X"E7",X"61",X"35",X"86",X"34",X"06",X"86",
		X"7F",X"97",X"04",X"1F",X"20",X"BD",X"F2",X"C3",X"BD",X"F3",X"54",X"35",X"86",X"34",X"06",X"86",
		X"7F",X"97",X"04",X"A6",X"A4",X"E6",X"22",X"BD",X"F2",X"C3",X"BD",X"F3",X"54",X"35",X"86",X"34",
		X"16",X"1F",X"20",X"BD",X"F2",X"FC",X"E6",X"61",X"BD",X"F4",X"0E",X"35",X"96",X"34",X"16",X"1F",
		X"21",X"BD",X"F2",X"F2",X"E6",X"61",X"AE",X"62",X"BD",X"F4",X"0E",X"35",X"96",X"34",X"56",X"86",
		X"7F",X"97",X"04",X"BD",X"F3",X"73",X"35",X"D6",X"34",X"56",X"1F",X"20",X"BD",X"F2",X"FC",X"BD",
		X"F4",X"95",X"35",X"B6",X"BD",X"F2",X"A9",X"CC",X"FC",X"38",X"FD",X"C8",X"2A",X"B6",X"C8",X"9B",
		X"10",X"8E",X"ED",X"A3",X"10",X"AE",X"A6",X"CE",X"ED",X"9F",X"EE",X"C6",X"8D",X"DA",X"39",X"BD",
		X"F2",X"A9",X"CC",X"FC",X"38",X"FD",X"C8",X"2A",X"10",X"8E",X"7F",X"A0",X"CE",X"C8",X"A8",X"8D",
		X"C7",X"B6",X"C8",X"79",X"27",X"09",X"10",X"8E",X"7F",X"10",X"CE",X"C8",X"AF",X"8D",X"B9",X"39",
		X"BD",X"F1",X"92",X"34",X"08",X"BD",X"F2",X"E6",X"BD",X"EA",X"B4",X"B6",X"C8",X"80",X"BD",X"F1",
		X"B4",X"FC",X"C8",X"81",X"FD",X"C8",X"1F",X"FD",X"C8",X"21",X"BD",X"F1",X"F8",X"86",X"C8",X"1F",
		X"8B",X"96",X"9C",X"27",X"08",X"0A",X"9C",X"26",X"04",X"AD",X"9F",X"C8",X"9D",X"96",X"9F",X"27",
		X"08",X"0A",X"9F",X"26",X"04",X"AD",X"9F",X"C8",X"A0",X"96",X"A2",X"27",X"08",X"0A",X"A2",X"26",
		X"04",X"AD",X"9F",X"C8",X"A3",X"96",X"A5",X"27",X"08",X"0A",X"A5",X"26",X"04",X"AD",X"9F",X"C8",
		X"A6",X"35",X"88",X"96",X"EA",X"27",X"12",X"10",X"8E",X"C9",X"0B",X"86",X"04",X"97",X"8F",X"6D",
		X"A4",X"26",X"07",X"31",X"2A",X"0A",X"8F",X"26",X"F6",X"39",X"96",X"E7",X"27",X"35",X"34",X"20",
		X"A6",X"25",X"E6",X"27",X"1F",X"01",X"CC",X"06",X"16",X"10",X"9E",X"DC",X"BD",X"F8",X"FF",X"35",
		X"20",X"24",X"20",X"6F",X"A4",X"0F",X"E7",X"0F",X"A2",X"8E",X"ED",X"9F",X"96",X"9B",X"AE",X"86",
		X"CC",X"10",X"00",X"BD",X"F8",X"7C",X"86",X"30",X"C6",X"70",X"9E",X"DC",X"BD",X"E7",X"84",X"0A",
		X"EA",X"20",X"C6",X"CE",X"C9",X"33",X"86",X"1C",X"97",X"90",X"A6",X"C4",X"84",X"3F",X"26",X"09",
		X"33",X"C8",X"12",X"0A",X"90",X"26",X"F3",X"20",X"AA",X"34",X"20",X"A6",X"25",X"E6",X"27",X"1F",
		X"01",X"A6",X"44",X"E6",X"46",X"1F",X"02",X"EC",X"4C",X"BD",X"F8",X"FF",X"35",X"20",X"24",X"E0",
		X"A6",X"41",X"84",X"02",X"27",X"5A",X"8E",X"ED",X"9F",X"96",X"9B",X"AE",X"86",X"EC",X"4E",X"BD",
		X"F8",X"7C",X"0C",X"F5",X"A6",X"44",X"E6",X"46",X"1F",X"01",X"A6",X"42",X"C6",X"20",X"BD",X"E7",
		X"84",X"CC",X"01",X"10",X"ED",X"4E",X"96",X"C8",X"A0",X"44",X"D6",X"CA",X"E0",X"46",X"BD",X"F5",
		X"93",X"80",X"10",X"1F",X"89",X"34",X"20",X"86",X"3F",X"BD",X"E7",X"B5",X"10",X"AF",X"48",X"AF",
		X"4A",X"35",X"20",X"6F",X"A4",X"CC",X"04",X"04",X"ED",X"4C",X"A6",X"41",X"E6",X"43",X"5A",X"27",
		X"06",X"BD",X"E9",X"A1",X"BD",X"E9",X"A1",X"86",X"04",X"A7",X"41",X"0A",X"EA",X"7E",X"EB",X"53",
		X"86",X"01",X"A7",X"C4",X"6F",X"A4",X"8E",X"ED",X"9F",X"96",X"9B",X"AE",X"86",X"EC",X"4E",X"BD",
		X"F8",X"7C",X"A6",X"44",X"E6",X"46",X"1F",X"01",X"A6",X"42",X"C6",X"40",X"BD",X"E7",X"84",X"0A",
		X"EB",X"0A",X"EA",X"7E",X"EB",X"53",X"96",X"BD",X"26",X"19",X"96",X"EE",X"26",X"15",X"10",X"8E",
		X"C9",X"33",X"86",X"1C",X"97",X"8F",X"A6",X"A4",X"84",X"3F",X"26",X"08",X"31",X"A8",X"12",X"0A",
		X"8F",X"26",X"F3",X"39",X"34",X"20",X"96",X"C8",X"D6",X"CA",X"1F",X"01",X"A6",X"24",X"E6",X"26",
		X"10",X"AE",X"2C",X"1E",X"20",X"BD",X"F8",X"FF",X"35",X"20",X"24",X"E0",X"6F",X"A4",X"0F",X"ED",
		X"96",X"C8",X"D6",X"CA",X"1F",X"01",X"A6",X"22",X"8A",X"80",X"C6",X"30",X"BD",X"E7",X"84",X"0C",
		X"F3",X"0A",X"EB",X"20",X"CE",X"96",X"BD",X"26",X"19",X"96",X"EE",X"26",X"15",X"96",X"E7",X"27",
		X"11",X"96",X"C8",X"D6",X"CA",X"1F",X"01",X"CC",X"06",X"16",X"10",X"9E",X"DC",X"BD",X"F8",X"FF",
		X"25",X"01",X"39",X"0F",X"E7",X"0F",X"A2",X"96",X"C8",X"D6",X"CA",X"1F",X"01",X"86",X"08",X"8A",
		X"80",X"C6",X"30",X"BD",X"E7",X"84",X"0C",X"F3",X"39",X"B6",X"C8",X"F2",X"27",X"08",X"7F",X"C8",
		X"F2",X"CE",X"ED",X"37",X"20",X"31",X"B6",X"C8",X"F3",X"27",X"08",X"7F",X"C8",X"F3",X"CE",X"ED",
		X"4D",X"20",X"24",X"B6",X"C8",X"B6",X"27",X"08",X"7F",X"C8",X"B6",X"CE",X"ED",X"42",X"20",X"17",
		X"B6",X"C8",X"F4",X"27",X"0B",X"7F",X"C8",X"F4",X"7F",X"C8",X"F6",X"CE",X"ED",X"5A",X"20",X"07",
		X"B6",X"C8",X"F6",X"26",X"F0",X"20",X"03",X"BD",X"F2",X"7D",X"F6",X"C8",X"00",X"CB",X"10",X"C1",
		X"A0",X"24",X"07",X"86",X"00",X"BD",X"F2",X"56",X"20",X"06",X"CC",X"08",X"00",X"BD",X"F2",X"56",
		X"F6",X"C8",X"02",X"CB",X"20",X"C1",X"F0",X"24",X"07",X"86",X"02",X"BD",X"F2",X"56",X"20",X"06",
		X"CC",X"09",X"00",X"BD",X"F2",X"56",X"39",X"00",X"10",X"01",X"00",X"06",X"1F",X"07",X"06",X"08",
		X"0F",X"FF",X"02",X"39",X"03",X"00",X"06",X"1F",X"07",X"05",X"09",X"0F",X"FF",X"06",X"1F",X"07",
		X"07",X"0A",X"10",X"0B",X"00",X"0C",X"38",X"0D",X"00",X"FF",X"00",X"00",X"01",X"00",X"02",X"30",
		X"03",X"00",X"04",X"00",X"05",X"00",X"06",X"1F",X"07",X"3D",X"08",X"00",X"09",X"0F",X"0A",X"00",
		X"0B",X"00",X"0C",X"00",X"0D",X"00",X"FF",X"ED",X"8F",X"FE",X"B6",X"00",X"19",X"01",X"19",X"00",
		X"19",X"01",X"32",X"00",X"19",X"01",X"19",X"00",X"19",X"06",X"19",X"05",X"19",X"00",X"80",X"FF",
		X"EE",X"DD",X"CC",X"BB",X"AA",X"99",X"88",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"C8",
		X"A8",X"C8",X"AF",X"7F",X"A0",X"7F",X"10",X"C8",X"F9",X"C9",X"00",X"86",X"0C",X"A0",X"84",X"A0",
		X"01",X"A0",X"02",X"A0",X"03",X"27",X"20",X"E6",X"84",X"CB",X"FD",X"C4",X"03",X"E7",X"84",X"C6",
		X"FC",X"E9",X"01",X"C4",X"03",X"E7",X"01",X"C6",X"FC",X"E9",X"02",X"C4",X"03",X"E7",X"02",X"C6",
		X"FC",X"E9",X"03",X"C4",X"03",X"E7",X"03",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C8",X"40",X"3F",X"00",X"20",X"80",X"10",X"1F",X"3F",X"3F",X"00",X"BF",X"BF",X"BF",X"C0",X"20",
		X"48",X"08",X"F8",X"30",X"A8",X"10",X"D0",X"A0",X"BF",X"BF",X"00",X"3F",X"3F",X"48",X"20",X"80",
		X"00",X"B0",X"48",X"38",X"FB",X"38",X"80",X"28",X"30",X"48",X"80",X"80",X"45",X"F0",X"28",X"7F",
		X"3F",X"BF",X"A5",X"00",X"D0",X"60",X"20",X"28",X"B8",X"40",X"15",X"80",X"40",X"F8",X"40",X"18",
		X"FA",X"38",X"E0",X"C0",X"4D",X"49",X"4E",X"45",X"20",X"46",X"49",X"45",X"4C",X"44",X"80",X"FA",
		X"38",X"E0",X"D8",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"80",X"00",X"10",X"00",
		X"FF",X"20",X"A0",X"FF",X"C0",X"40",X"FF",X"90",X"20",X"FF",X"70",X"20",X"FF",X"50",X"50",X"FF",
		X"D0",X"90",X"01",X"00",X"20",X"00",X"FF",X"30",X"B0",X"FF",X"B0",X"30",X"FF",X"B0",X"D0",X"FF",
		X"30",X"50",X"FF",X"D0",X"50",X"FF",X"50",X"D0",X"FF",X"50",X"30",X"FF",X"D0",X"B0",X"01",X"FF",
		X"00",X"00",X"00",X"30",X"00",X"FF",X"10",X"C0",X"FF",X"C0",X"10",X"FF",X"C0",X"F0",X"FF",X"10",
		X"40",X"FF",X"F0",X"40",X"FF",X"40",X"F0",X"FF",X"40",X"10",X"FF",X"F0",X"C0",X"01",X"FF",X"00",
		X"00",X"00",X"F0",X"D0",X"FF",X"C0",X"40",X"FF",X"20",X"00",X"FF",X"40",X"40",X"FF",X"00",X"E0",
		X"FF",X"40",X"C0",X"FF",X"E0",X"00",X"FF",X"C0",X"C0",X"FF",X"00",X"20",X"01",X"00",X"3F",X"00",
		X"FF",X"80",X"00",X"00",X"3F",X"3F",X"FF",X"00",X"80",X"01",X"FF",X"7F",X"20",X"00",X"C0",X"10",
		X"FF",X"C0",X"D0",X"FF",X"20",X"7F",X"00",X"E0",X"C0",X"FF",X"00",X"C0",X"FF",X"E0",X"30",X"00",
		X"C0",X"00",X"FF",X"60",X"CD",X"FF",X"A0",X"00",X"00",X"20",X"D0",X"FF",X"3C",X"30",X"FF",X"00",
		X"82",X"00",X"30",X"30",X"FF",X"D0",X"50",X"FF",X"20",X"F0",X"01",X"00",X"3F",X"00",X"FF",X"C4",
		X"08",X"FF",X"D8",X"D8",X"FF",X"20",X"00",X"00",X"00",X"40",X"FF",X"E0",X"00",X"FF",X"28",X"D8",
		X"FF",X"3C",X"08",X"01",X"00",X"3F",X"00",X"FF",X"C4",X"08",X"01",X"00",X"04",X"08",X"FF",X"D8",
		X"D8",X"FF",X"20",X"00",X"01",X"00",X"3F",X"00",X"FF",X"C4",X"F8",X"01",X"00",X"04",X"F8",X"FF",
		X"D8",X"28",X"FF",X"20",X"00",X"01",X"00",X"20",X"00",X"FF",X"00",X"D8",X"FF",X"D0",X"A8",X"FF",
		X"F0",X"40",X"FF",X"08",X"18",X"FF",X"18",X"F0",X"FF",X"F0",X"B8",X"00",X"10",X"48",X"FF",X"08",
		X"00",X"FF",X"E8",X"10",X"FF",X"F8",X"00",X"00",X"08",X"00",X"FF",X"00",X"06",X"00",X"10",X"FA",
		X"FF",X"08",X"00",X"FF",X"00",X"F0",X"00",X"10",X"18",X"FF",X"F0",X"08",X"01",X"00",X"20",X"00",
		X"FF",X"00",X"28",X"FF",X"D0",X"58",X"FF",X"F0",X"C0",X"FF",X"08",X"E8",X"FF",X"18",X"10",X"FF",
		X"F0",X"48",X"00",X"10",X"B8",X"FF",X"08",X"00",X"FF",X"E8",X"F0",X"FF",X"F8",X"00",X"FF",X"08",
		X"00",X"FF",X"00",X"FA",X"00",X"10",X"06",X"FF",X"08",X"00",X"FF",X"00",X"10",X"00",X"10",X"E8",
		X"FF",X"F0",X"F8",X"01",X"FF",X"00",X"D8",X"FF",X"E8",X"08",X"FF",X"00",X"40",X"FF",X"18",X"08",
		X"FF",X"00",X"D8",X"00",X"08",X"E0",X"FF",X"10",X"00",X"FF",X"00",X"40",X"FF",X"F0",X"00",X"FF",
		X"00",X"C0",X"01",X"00",X"18",X"00",X"FF",X"00",X"20",X"FF",X"C8",X"70",X"FF",X"10",X"A0",X"FF",
		X"00",X"A0",X"FF",X"EC",X"A4",X"FF",X"39",X"6D",X"FF",X"00",X"20",X"01",X"7F",X"C8",X"25",X"7F",
		X"C8",X"26",X"7F",X"C8",X"3B",X"7E",X"F0",X"1C",X"B6",X"C8",X"D9",X"27",X"09",X"81",X"08",X"2F",
		X"02",X"86",X"08",X"B7",X"C8",X"8F",X"39",X"BD",X"F1",X"BA",X"BD",X"F1",X"AF",X"96",X"0F",X"10",
		X"26",X"00",X"79",X"7E",X"F0",X"1F",X"67",X"20",X"4D",X"42",X"20",X"80",X"00",X"00",X"00",X"00",
		X"10",X"CE",X"CB",X"EA",X"BD",X"F1",X"8B",X"CC",X"73",X"21",X"10",X"B3",X"CB",X"FE",X"27",X"5C",
		X"FD",X"CB",X"FE",X"7C",X"C8",X"3B",X"8E",X"CB",X"EB",X"BD",X"F8",X"4F",X"BD",X"F1",X"AF",X"DC",
		X"25",X"10",X"83",X"01",X"01",X"26",X"02",X"D7",X"56",X"57",X"C4",X"03",X"8E",X"F0",X"FD",X"E6",
		X"85",X"D7",X"29",X"C6",X"02",X"D7",X"24",X"CE",X"FD",X"0D",X"BD",X"F6",X"87",X"BD",X"F1",X"92",
		X"BD",X"F2",X"89",X"BD",X"F2",X"A9",X"B6",X"C8",X"26",X"CE",X"F1",X"0C",X"85",X"20",X"27",X"02",
		X"33",X"4C",X"BD",X"F3",X"85",X"8E",X"F0",X"E9",X"BD",X"F3",X"08",X"86",X"03",X"BD",X"F4",X"34",
		X"7A",X"C8",X"24",X"26",X"F3",X"B6",X"C8",X"25",X"81",X"01",X"23",X"B0",X"BD",X"F1",X"AF",X"86",
		X"CC",X"97",X"29",X"CC",X"F1",X"01",X"DD",X"39",X"0F",X"25",X"0F",X"26",X"CE",X"00",X"00",X"8E",
		X"F1",X"01",X"C6",X"0B",X"A6",X"C0",X"A1",X"80",X"27",X"0D",X"C1",X"01",X"27",X"04",X"C1",X"05",
		X"23",X"05",X"CE",X"E0",X"00",X"20",X"07",X"5A",X"26",X"EA",X"D7",X"39",X"D7",X"3A",X"0C",X"56",
		X"DF",X"37",X"EE",X"C4",X"BD",X"F1",X"AF",X"CC",X"F8",X"48",X"DD",X"2A",X"BD",X"F6",X"87",X"BD",
		X"F1",X"92",X"BD",X"F2",X"89",X"BD",X"F2",X"A9",X"CC",X"C0",X"C0",X"FE",X"C8",X"39",X"BD",X"F3",
		X"7A",X"B6",X"C8",X"3B",X"26",X"0C",X"4A",X"CE",X"CB",X"EB",X"A7",X"46",X"CC",X"68",X"D0",X"BD",
		X"F3",X"7A",X"FE",X"C8",X"37",X"33",X"42",X"BD",X"F3",X"85",X"B6",X"C8",X"56",X"26",X"C5",X"BE",
		X"C8",X"25",X"8C",X"00",X"7D",X"23",X"BD",X"6E",X"41",X"40",X"D6",X"00",X"56",X"81",X"00",X"00",
		X"A9",X"7E",X"00",X"39",X"DC",X"8E",X"00",X"00",X"4A",X"72",X"00",X"00",X"B6",X"E0",X"38",X"0E",
		X"03",X"67",X"20",X"47",X"43",X"45",X"20",X"31",X"39",X"38",X"32",X"80",X"F1",X"60",X"27",X"CF",
		X"56",X"45",X"43",X"54",X"52",X"45",X"58",X"80",X"F3",X"60",X"26",X"CF",X"56",X"45",X"43",X"54",
		X"52",X"45",X"58",X"80",X"FC",X"60",X"DF",X"E9",X"47",X"43",X"45",X"80",X"FC",X"38",X"CC",X"D1",
		X"45",X"4E",X"54",X"45",X"52",X"54",X"41",X"49",X"4E",X"49",X"4E",X"47",X"80",X"FC",X"38",X"BC",
		X"DC",X"4E",X"45",X"57",X"20",X"49",X"44",X"45",X"41",X"53",X"80",X"00",X"8D",X"5C",X"CC",X"9F",
		X"FF",X"DD",X"02",X"CC",X"01",X"00",X"DD",X"00",X"CC",X"98",X"7F",X"97",X"0B",X"D7",X"04",X"BD",
		X"F3",X"54",X"20",X"3E",X"8D",X"49",X"C6",X"7A",X"8E",X"C8",X"00",X"BD",X"F5",X"3F",X"CC",X"C8",
		X"7D",X"DD",X"7B",X"0C",X"7D",X"27",X"FC",X"86",X"05",X"97",X"28",X"CC",X"30",X"75",X"DD",X"3D",
		X"CC",X"01",X"03",X"DD",X"1F",X"CC",X"05",X"07",X"DD",X"21",X"39",X"8D",X"D7",X"8D",X"BD",X"7E",
		X"F2",X"72",X"BE",X"C8",X"25",X"30",X"01",X"BF",X"C8",X"25",X"8D",X"0E",X"86",X"20",X"95",X"0D",
		X"27",X"FC",X"FC",X"C8",X"3D",X"DD",X"08",X"7E",X"F2",X"E6",X"86",X"D0",X"1F",X"8B",X"39",X"86",
		X"C8",X"1F",X"8B",X"39",X"B4",X"C8",X"0F",X"B7",X"C8",X"0F",X"8E",X"C8",X"12",X"A6",X"1D",X"A7",
		X"1E",X"86",X"0E",X"97",X"01",X"CC",X"19",X"01",X"97",X"00",X"12",X"D7",X"00",X"0F",X"03",X"CC",
		X"09",X"01",X"97",X"00",X"12",X"96",X"01",X"43",X"A7",X"1D",X"D7",X"00",X"C6",X"FF",X"D7",X"03",
		X"43",X"AA",X"1E",X"43",X"A7",X"1F",X"34",X"02",X"C6",X"01",X"1F",X"98",X"A4",X"E4",X"A7",X"80",
		X"58",X"26",X"F7",X"35",X"82",X"7A",X"C8",X"23",X"8E",X"C8",X"1F",X"A6",X"80",X"26",X"0C",X"8C",
		X"C8",X"23",X"26",X"F7",X"6F",X"84",X"86",X"01",X"97",X"00",X"39",X"97",X"00",X"0F",X"01",X"0A",
		X"00",X"C6",X"60",X"5C",X"2A",X"FD",X"B6",X"C8",X"23",X"2B",X"25",X"86",X"20",X"0C",X"00",X"95",
		X"00",X"27",X"0A",X"C6",X"40",X"D7",X"01",X"95",X"00",X"26",X"0B",X"20",X"08",X"C6",X"C0",X"D7",
		X"01",X"95",X"00",X"27",X"01",X"5F",X"E7",X"1B",X"20",X"C5",X"1F",X"98",X"9A",X"01",X"97",X"01",
		X"86",X"20",X"95",X"00",X"26",X"06",X"1F",X"98",X"98",X"01",X"97",X"01",X"54",X"F1",X"C8",X"1A",
		X"26",X"E8",X"D6",X"01",X"20",X"E0",X"8E",X"C8",X"00",X"E7",X"86",X"97",X"01",X"86",X"19",X"97",
		X"00",X"86",X"01",X"97",X"00",X"96",X"01",X"D7",X"01",X"C6",X"11",X"D7",X"00",X"C6",X"01",X"D7",
		X"00",X"39",X"CC",X"0E",X"00",X"8D",X"DF",X"4A",X"2A",X"FB",X"7E",X"F5",X"33",X"8E",X"C8",X"00",
		X"20",X"02",X"8D",X"D5",X"EC",X"C1",X"2A",X"FA",X"39",X"8E",X"C8",X"00",X"CE",X"C8",X"3F",X"86",
		X"0D",X"E6",X"C0",X"E1",X"86",X"27",X"02",X"8D",X"C0",X"4A",X"2A",X"F5",X"39",X"86",X"1F",X"20",
		X"0A",X"86",X"3F",X"20",X"06",X"86",X"5F",X"20",X"02",X"86",X"7F",X"97",X"01",X"B7",X"C8",X"27",
		X"CC",X"05",X"04",X"97",X"00",X"D7",X"00",X"D7",X"00",X"C6",X"01",X"D7",X"00",X"39",X"F7",X"C8",
		X"28",X"EC",X"81",X"8D",X"4D",X"86",X"FF",X"97",X"0A",X"F6",X"C8",X"28",X"5A",X"26",X"FD",X"0F",
		X"0A",X"39",X"7A",X"C8",X"23",X"8D",X"EA",X"B6",X"C8",X"23",X"26",X"F6",X"20",X"76",X"A6",X"80",
		X"2E",X"72",X"8D",X"DD",X"20",X"F8",X"8E",X"F9",X"F0",X"8D",X"1D",X"BD",X"F3",X"6B",X"8D",X"20",
		X"20",X"62",X"C6",X"7F",X"D7",X"04",X"A6",X"84",X"E6",X"02",X"20",X"16",X"97",X"01",X"34",X"06",
		X"86",X"7F",X"97",X"04",X"0F",X"00",X"20",X"10",X"C6",X"FF",X"20",X"02",X"C6",X"7F",X"D7",X"04",
		X"EC",X"81",X"97",X"01",X"0F",X"00",X"34",X"06",X"86",X"CE",X"97",X"0C",X"0F",X"0A",X"0C",X"00",
		X"D7",X"01",X"0F",X"05",X"35",X"06",X"BD",X"F5",X"84",X"E7",X"7F",X"AA",X"7F",X"C6",X"40",X"81",
		X"40",X"23",X"12",X"81",X"64",X"23",X"04",X"86",X"08",X"20",X"02",X"86",X"04",X"D5",X"0D",X"27",
		X"FC",X"4A",X"26",X"FD",X"39",X"D5",X"0D",X"27",X"FC",X"39",X"BD",X"F1",X"AA",X"20",X"05",X"B6",
		X"C8",X"24",X"27",X"16",X"CC",X"00",X"CC",X"D7",X"0C",X"97",X"0A",X"CC",X"03",X"02",X"0F",X"01",
		X"97",X"00",X"D7",X"00",X"D7",X"00",X"C6",X"01",X"D7",X"00",X"39",X"CC",X"00",X"CC",X"D7",X"0C",
		X"97",X"0A",X"39",X"EC",X"C1",X"FD",X"C8",X"2A",X"EC",X"C1",X"BD",X"F2",X"FC",X"BD",X"F5",X"75",
		X"7E",X"F4",X"95",X"8D",X"EE",X"A6",X"C4",X"26",X"FA",X"39",X"8D",X"EC",X"A6",X"C4",X"26",X"FA",
		X"39",X"AE",X"84",X"34",X"04",X"C6",X"80",X"33",X"78",X"36",X"06",X"35",X"02",X"81",X"09",X"23",
		X"02",X"86",X"3C",X"8B",X"30",X"C6",X"2D",X"36",X"06",X"36",X"10",X"20",X"CB",X"A6",X"80",X"20",
		X"08",X"D7",X"04",X"20",X"07",X"EC",X"81",X"D7",X"04",X"B7",X"C8",X"23",X"EC",X"84",X"97",X"01",
		X"0F",X"00",X"30",X"02",X"12",X"0C",X"00",X"D7",X"01",X"CC",X"00",X"00",X"20",X"1F",X"A6",X"80",
		X"20",X"08",X"D7",X"04",X"20",X"07",X"EC",X"81",X"D7",X"04",X"B7",X"C8",X"23",X"EC",X"84",X"97",
		X"01",X"0F",X"00",X"30",X"02",X"12",X"0C",X"00",X"D7",X"01",X"CC",X"FF",X"00",X"97",X"0A",X"D7",
		X"05",X"CC",X"00",X"40",X"D5",X"0D",X"27",X"FC",X"12",X"97",X"0A",X"B6",X"C8",X"23",X"4A",X"2A",
		X"D9",X"7E",X"F3",X"4F",X"C6",X"FF",X"20",X"06",X"C6",X"7F",X"20",X"02",X"E6",X"80",X"D7",X"04",
		X"EC",X"01",X"97",X"01",X"0F",X"00",X"A6",X"84",X"30",X"03",X"0C",X"00",X"D7",X"01",X"97",X"0A",
		X"0F",X"05",X"CC",X"00",X"40",X"D5",X"0D",X"27",X"FC",X"12",X"97",X"0A",X"A6",X"84",X"2F",X"E0",
		X"7E",X"F3",X"4F",X"4A",X"B7",X"C8",X"23",X"EC",X"84",X"97",X"01",X"0F",X"00",X"30",X"02",X"0C",
		X"00",X"D7",X"01",X"B6",X"C8",X"29",X"C6",X"40",X"97",X"0A",X"0F",X"05",X"F5",X"D0",X"0D",X"27",
		X"0B",X"0F",X"0A",X"B6",X"C8",X"23",X"26",X"DB",X"39",X"B6",X"C8",X"29",X"97",X"0A",X"12",X"D5",
		X"0D",X"27",X"F6",X"B6",X"C8",X"23",X"0F",X"0A",X"4D",X"26",X"C8",X"7E",X"F3",X"4F",X"B6",X"C8",
		X"24",X"34",X"02",X"7F",X"C8",X"24",X"A6",X"80",X"2A",X"04",X"8D",X"BB",X"20",X"F8",X"26",X"05",
		X"BD",X"F3",X"BC",X"20",X"F1",X"4A",X"27",X"05",X"BD",X"F3",X"DD",X"20",X"E9",X"35",X"02",X"B7",
		X"C8",X"24",X"7E",X"F3",X"4F",X"FF",X"C8",X"2C",X"8E",X"F9",X"D4",X"CC",X"18",X"83",X"0F",X"01",
		X"97",X"0B",X"8E",X"F9",X"D4",X"D7",X"00",X"0A",X"00",X"CC",X"80",X"81",X"12",X"0C",X"00",X"D7",
		X"00",X"97",X"00",X"7D",X"C8",X"00",X"0C",X"00",X"B6",X"C8",X"2B",X"97",X"01",X"CC",X"01",X"00",
		X"FE",X"C8",X"2C",X"97",X"00",X"20",X"04",X"A6",X"86",X"97",X"0A",X"A6",X"C0",X"2A",X"F8",X"86",
		X"81",X"97",X"00",X"00",X"01",X"86",X"01",X"97",X"00",X"8C",X"FB",X"B4",X"27",X"2C",X"30",X"88",
		X"50",X"1F",X"30",X"B3",X"C8",X"2C",X"C0",X"02",X"58",X"21",X"00",X"86",X"81",X"12",X"5A",X"26",
		X"FA",X"97",X"00",X"F6",X"C8",X"2A",X"D7",X"01",X"0A",X"00",X"CC",X"81",X"01",X"12",X"97",X"00",
		X"0F",X"01",X"D7",X"00",X"97",X"00",X"C6",X"03",X"20",X"9B",X"86",X"98",X"97",X"0B",X"7E",X"F3",
		X"54",X"34",X"14",X"C6",X"02",X"20",X"03",X"34",X"14",X"5F",X"BE",X"C8",X"7B",X"A6",X"01",X"49",
		X"49",X"49",X"49",X"A8",X"02",X"46",X"69",X"84",X"69",X"01",X"69",X"02",X"5A",X"2A",X"EE",X"A6",
		X"84",X"35",X"94",X"C6",X"0D",X"8E",X"C8",X"3F",X"8D",X"05",X"86",X"3F",X"A7",X"06",X"39",X"4F",
		X"20",X"06",X"8E",X"C8",X"00",X"CC",X"00",X"FF",X"6F",X"8B",X"83",X"00",X"01",X"2A",X"F9",X"39",
		X"86",X"80",X"A7",X"85",X"5A",X"26",X"FB",X"A7",X"84",X"39",X"C6",X"02",X"20",X"02",X"C6",X"05",
		X"8E",X"C8",X"2E",X"6D",X"85",X"27",X"02",X"6A",X"85",X"5A",X"2A",X"F7",X"39",X"C6",X"03",X"20",
		X"09",X"C6",X"02",X"20",X"05",X"C6",X"01",X"20",X"01",X"5F",X"5A",X"2A",X"FD",X"39",X"8E",X"F9",
		X"DC",X"A6",X"86",X"39",X"4D",X"2A",X"04",X"40",X"28",X"01",X"4A",X"5D",X"2A",X"04",X"50",X"28",
		X"01",X"5A",X"39",X"34",X"10",X"DD",X"34",X"59",X"C6",X"00",X"59",X"49",X"59",X"58",X"D7",X"36",
		X"DC",X"34",X"8D",X"E0",X"97",X"34",X"D1",X"34",X"23",X"08",X"0C",X"36",X"1E",X"89",X"20",X"02",
		X"44",X"54",X"81",X"09",X"22",X"FA",X"DD",X"34",X"D6",X"36",X"8E",X"FC",X"24",X"E6",X"85",X"8E",
		X"FC",X"2C",X"A6",X"86",X"9B",X"35",X"8B",X"0A",X"C5",X"01",X"26",X"04",X"EB",X"86",X"20",X"03",
		X"5A",X"E0",X"86",X"D7",X"36",X"96",X"36",X"35",X"90",X"8B",X"10",X"8E",X"FC",X"6D",X"5F",X"85",
		X"20",X"27",X"02",X"C6",X"80",X"84",X"1F",X"81",X"10",X"26",X"01",X"5C",X"A6",X"86",X"39",X"34",
		X"10",X"96",X"36",X"8D",X"E6",X"DD",X"37",X"96",X"36",X"8D",X"DE",X"DD",X"39",X"35",X"90",X"C0",
		X"10",X"D7",X"36",X"97",X"3B",X"8D",X"E8",X"8D",X"54",X"40",X"34",X"02",X"8D",X"55",X"35",X"84",
		X"B7",X"C8",X"36",X"F7",X"C8",X"23",X"34",X"08",X"BD",X"F1",X"AF",X"8D",X"D2",X"20",X"18",X"B7",
		X"C8",X"36",X"34",X"08",X"BD",X"F1",X"AF",X"97",X"23",X"8D",X"C4",X"A6",X"80",X"A7",X"C0",X"2F",
		X"06",X"0F",X"23",X"35",X"88",X"0A",X"23",X"A6",X"80",X"8D",X"26",X"A7",X"C4",X"A6",X"84",X"8D",
		X"1A",X"AB",X"C4",X"A7",X"C0",X"A6",X"1F",X"8D",X"12",X"A7",X"C4",X"A6",X"80",X"8D",X"12",X"A0",
		X"C4",X"A7",X"C0",X"96",X"23",X"2B",X"D4",X"26",X"DC",X"35",X"88",X"97",X"3B",X"DC",X"37",X"20",
		X"04",X"97",X"3B",X"DC",X"39",X"D7",X"3C",X"C5",X"01",X"27",X"04",X"96",X"3B",X"20",X"0A",X"D6",
		X"3B",X"2A",X"03",X"03",X"3C",X"50",X"3D",X"89",X"00",X"D6",X"3C",X"2A",X"01",X"40",X"39",X"E6",
		X"C6",X"E7",X"86",X"4A",X"2A",X"F9",X"39",X"96",X"56",X"2B",X"28",X"27",X"F9",X"8E",X"FC",X"8D",
		X"9F",X"4D",X"86",X"80",X"97",X"56",X"EC",X"C1",X"DD",X"4F",X"EC",X"C1",X"DD",X"51",X"DF",X"53",
		X"BD",X"F5",X"33",X"CC",X"1F",X"1F",X"DD",X"5F",X"CC",X"00",X"00",X"DD",X"63",X"DD",X"65",X"97",
		X"55",X"20",X"39",X"CE",X"C8",X"5E",X"C6",X"02",X"A6",X"C5",X"81",X"1F",X"27",X"02",X"6C",X"C5",
		X"5A",X"2A",X"F5",X"9E",X"51",X"CE",X"C8",X"58",X"86",X"07",X"6C",X"C4",X"A1",X"C4",X"2C",X"02",
		X"6F",X"C4",X"E6",X"C0",X"C4",X"07",X"E6",X"85",X"E7",X"C0",X"4C",X"81",X"09",X"23",X"EB",X"0A",
		X"57",X"26",X"6B",X"96",X"55",X"4A",X"2A",X"02",X"86",X"02",X"97",X"55",X"E6",X"9F",X"C8",X"53",
		X"CE",X"C8",X"5E",X"6F",X"C6",X"C5",X"40",X"27",X"19",X"8E",X"F9",X"E4",X"A6",X"86",X"94",X"45",
		X"97",X"45",X"96",X"55",X"8B",X"03",X"A6",X"86",X"9A",X"45",X"97",X"45",X"C4",X"1F",X"D7",X"46",
		X"20",X"23",X"8E",X"F9",X"EA",X"A6",X"86",X"94",X"45",X"97",X"45",X"96",X"55",X"8B",X"03",X"A6",
		X"86",X"9A",X"45",X"97",X"45",X"96",X"55",X"48",X"8B",X"03",X"33",X"C6",X"C4",X"3F",X"58",X"9E",
		X"4D",X"EC",X"85",X"ED",X"C4",X"9E",X"53",X"E6",X"80",X"9F",X"53",X"5D",X"2B",X"A5",X"E6",X"80",
		X"2A",X"06",X"BD",X"F5",X"33",X"0F",X"56",X"39",X"9F",X"53",X"C4",X"3F",X"D7",X"57",X"10",X"9E",
		X"4F",X"CE",X"C8",X"5E",X"8E",X"C8",X"42",X"86",X"02",X"E6",X"C0",X"C5",X"01",X"27",X"07",X"54",
		X"E6",X"A5",X"C4",X"0F",X"20",X"07",X"54",X"E6",X"A5",X"54",X"54",X"54",X"54",X"E7",X"86",X"4A",
		X"2A",X"E7",X"CE",X"C8",X"67",X"8E",X"C8",X"47",X"EC",X"C3",X"6D",X"58",X"2A",X"0A",X"60",X"58",
		X"E0",X"58",X"82",X"00",X"60",X"58",X"20",X"04",X"EB",X"58",X"89",X"00",X"ED",X"81",X"8C",X"C8",
		X"4D",X"26",X"E5",X"39",X"20",X"C0",X"40",X"C0",X"50",X"4C",X"41",X"59",X"45",X"52",X"80",X"E0",
		X"C0",X"01",X"C0",X"20",X"47",X"41",X"4D",X"45",X"80",X"FD",X"C8",X"4F",X"4D",X"27",X"02",X"86",
		X"01",X"5D",X"27",X"02",X"C6",X"01",X"FD",X"C8",X"79",X"BD",X"F1",X"AF",X"CC",X"F8",X"50",X"DD",
		X"2A",X"97",X"3C",X"20",X"67",X"BD",X"F1",X"92",X"4F",X"BD",X"F1",X"B4",X"BD",X"F5",X"5A",X"BD",
		X"F2",X"A9",X"B6",X"C8",X"79",X"10",X"8E",X"F7",X"94",X"8D",X"5A",X"B6",X"C8",X"7A",X"10",X"8E",
		X"F7",X"9F",X"8D",X"51",X"BD",X"F1",X"AF",X"96",X"3C",X"27",X"06",X"96",X"0F",X"26",X"3D",X"0F",
		X"3C",X"96",X"2F",X"27",X"9E",X"96",X"2E",X"26",X"CC",X"96",X"15",X"26",X"96",X"96",X"12",X"27",
		X"0F",X"96",X"79",X"27",X"0B",X"4C",X"91",X"4F",X"23",X"02",X"86",X"01",X"97",X"79",X"20",X"1C",
		X"96",X"7A",X"27",X"B1",X"D6",X"13",X"27",X"09",X"4C",X"91",X"50",X"23",X"0D",X"86",X"01",X"20",
		X"09",X"D6",X"14",X"27",X"A0",X"4A",X"26",X"02",X"96",X"50",X"97",X"7A",X"86",X"F3",X"97",X"2F",
		X"43",X"97",X"2E",X"20",X"90",X"8E",X"C8",X"5E",X"34",X"02",X"8D",X"13",X"A6",X"E0",X"27",X"0E",
		X"8D",X"1C",X"1F",X"13",X"EC",X"A1",X"BD",X"F3",X"7A",X"1F",X"23",X"BD",X"F3",X"78",X"39",X"CC",
		X"20",X"20",X"ED",X"84",X"ED",X"02",X"A7",X"04",X"CC",X"30",X"80",X"ED",X"05",X"39",X"CE",X"00",
		X"00",X"81",X"63",X"23",X"08",X"80",X"64",X"33",X"C9",X"01",X"00",X"20",X"F4",X"81",X"09",X"23",
		X"07",X"80",X"0A",X"33",X"C8",X"10",X"20",X"F5",X"33",X"C6",X"1F",X"30",X"34",X"02",X"34",X"04",
		X"C6",X"05",X"4F",X"C1",X"01",X"23",X"10",X"C5",X"01",X"27",X"04",X"A6",X"E4",X"20",X"06",X"A6",
		X"E0",X"44",X"44",X"44",X"44",X"84",X"0F",X"BB",X"C8",X"23",X"7F",X"C8",X"23",X"AB",X"85",X"81",
		X"2F",X"2E",X"02",X"8B",X"10",X"81",X"39",X"23",X"05",X"80",X"0A",X"7C",X"C8",X"23",X"A7",X"85",
		X"5A",X"2A",X"CF",X"7F",X"C8",X"23",X"5F",X"A6",X"85",X"81",X"30",X"26",X"09",X"86",X"20",X"A7",
		X"85",X"5C",X"C1",X"05",X"2D",X"F1",X"39",X"34",X"50",X"4F",X"E6",X"80",X"2B",X"08",X"E1",X"C0",
		X"27",X"F8",X"22",X"01",X"4C",X"4C",X"35",X"D0",X"8D",X"ED",X"81",X"01",X"26",X"06",X"A6",X"80",
		X"A7",X"C0",X"2A",X"FA",X"39",X"34",X"20",X"34",X"36",X"EC",X"64",X"AB",X"C4",X"EB",X"41",X"ED",
		X"64",X"20",X"10",X"34",X"20",X"34",X"36",X"1F",X"30",X"AB",X"64",X"EB",X"65",X"20",X"F0",X"34",
		X"20",X"34",X"36",X"1F",X"41",X"5F",X"3A",X"A6",X"04",X"AB",X"84",X"28",X"02",X"86",X"7F",X"A1",
		X"02",X"2D",X"15",X"A6",X"04",X"A0",X"84",X"28",X"02",X"86",X"80",X"A1",X"02",X"2E",X"09",X"5C",
		X"C1",X"02",X"25",X"E2",X"1A",X"01",X"20",X"02",X"1C",X"FE",X"35",X"36",X"35",X"A0",X"96",X"67",
		X"2A",X"29",X"84",X"7F",X"97",X"67",X"8E",X"C8",X"58",X"86",X"04",X"BD",X"F6",X"83",X"54",X"54",
		X"54",X"DA",X"58",X"C4",X"07",X"D7",X"54",X"D6",X"58",X"C4",X"38",X"D7",X"53",X"D6",X"58",X"C4",
		X"07",X"D7",X"5D",X"C6",X"02",X"D7",X"5C",X"86",X"7F",X"20",X"0D",X"96",X"77",X"27",X"6A",X"90",
		X"5B",X"2A",X"05",X"5F",X"D7",X"77",X"20",X"62",X"97",X"77",X"44",X"44",X"D6",X"53",X"27",X"0D",
		X"97",X"46",X"D6",X"59",X"2B",X"05",X"27",X"05",X"1F",X"89",X"53",X"D7",X"46",X"44",X"81",X"07",
		X"23",X"05",X"81",X"0F",X"27",X"01",X"4C",X"D6",X"5A",X"2B",X"06",X"27",X"02",X"88",X"0F",X"1F",
		X"89",X"8D",X"37",X"D6",X"5D",X"27",X"2B",X"96",X"5C",X"4A",X"2A",X"02",X"86",X"02",X"97",X"5C",
		X"BD",X"F5",X"7E",X"95",X"5D",X"27",X"F0",X"D6",X"5C",X"58",X"50",X"8E",X"C8",X"4B",X"30",X"85",
		X"BD",X"F5",X"17",X"84",X"0F",X"81",X"05",X"22",X"03",X"48",X"8B",X"05",X"A7",X"84",X"96",X"7E",
		X"A7",X"01",X"96",X"58",X"43",X"94",X"45",X"97",X"45",X"39",X"96",X"54",X"8E",X"C8",X"45",X"4D",
		X"27",X"09",X"30",X"1F",X"44",X"24",X"F8",X"E7",X"84",X"20",X"F4",X"39",X"01",X"02",X"04",X"08",
		X"10",X"20",X"40",X"80",X"F7",X"EF",X"DF",X"01",X"02",X"04",X"FE",X"FD",X"FB",X"08",X"10",X"20",
		X"7F",X"7F",X"80",X"80",X"00",X"20",X"50",X"50",X"20",X"C8",X"20",X"10",X"10",X"40",X"20",X"00",
		X"00",X"00",X"00",X"08",X"30",X"20",X"70",X"70",X"10",X"F8",X"30",X"F8",X"70",X"70",X"00",X"60",
		X"00",X"00",X"00",X"70",X"70",X"20",X"F0",X"70",X"F0",X"F8",X"F8",X"78",X"88",X"70",X"08",X"88",
		X"80",X"88",X"88",X"F8",X"F0",X"70",X"F0",X"70",X"F8",X"88",X"88",X"88",X"88",X"88",X"F8",X"70",
		X"80",X"70",X"20",X"00",X"00",X"20",X"08",X"20",X"00",X"00",X"00",X"38",X"10",X"20",X"44",X"44",
		X"00",X"FE",X"FF",X"FE",X"00",X"70",X"50",X"50",X"78",X"C8",X"50",X"20",X"20",X"20",X"A8",X"20",
		X"00",X"00",X"00",X"08",X"48",X"60",X"88",X"88",X"30",X"80",X"40",X"08",X"88",X"88",X"60",X"60",
		X"10",X"00",X"40",X"88",X"88",X"50",X"48",X"88",X"48",X"80",X"80",X"80",X"88",X"20",X"08",X"90",
		X"80",X"D8",X"C8",X"88",X"88",X"88",X"88",X"88",X"A8",X"88",X"88",X"88",X"88",X"88",X"08",X"40",
		X"80",X"08",X"50",X"00",X"00",X"70",X"0C",X"20",X"70",X"70",X"00",X"44",X"10",X"70",X"00",X"00",
		X"6C",X"82",X"FF",X"FE",X"00",X"70",X"50",X"F8",X"A0",X"10",X"50",X"40",X"40",X"10",X"70",X"20",
		X"00",X"00",X"00",X"10",X"48",X"20",X"08",X"08",X"50",X"F0",X"80",X"10",X"88",X"88",X"60",X"00",
		X"20",X"78",X"20",X"08",X"A8",X"88",X"48",X"80",X"48",X"80",X"80",X"80",X"88",X"20",X"08",X"A0",
		X"80",X"A8",X"A8",X"88",X"88",X"88",X"88",X"40",X"20",X"88",X"88",X"88",X"50",X"50",X"10",X"40",
		X"40",X"08",X"88",X"00",X"70",X"A8",X"0A",X"20",X"88",X"F8",X"60",X"BA",X"38",X"20",X"00",X"00",
		X"92",X"82",X"FF",X"FE",X"00",X"20",X"00",X"50",X"70",X"20",X"60",X"00",X"40",X"10",X"A8",X"F8",
		X"00",X"70",X"00",X"20",X"48",X"20",X"70",X"30",X"90",X"08",X"F0",X"20",X"70",X"78",X"00",X"60",
		X"40",X"00",X"10",X"10",X"B8",X"88",X"70",X"80",X"48",X"E0",X"E0",X"98",X"F8",X"20",X"08",X"C0",
		X"80",X"A8",X"98",X"88",X"F0",X"88",X"F0",X"20",X"20",X"88",X"50",X"A8",X"20",X"20",X"20",X"40",
		X"20",X"08",X"00",X"00",X"FE",X"20",X"08",X"20",X"88",X"F8",X"F0",X"A2",X"38",X"F8",X"82",X"38",
		X"92",X"82",X"FF",X"FE",X"00",X"00",X"00",X"F8",X"70",X"40",X"A8",X"00",X"40",X"10",X"A8",X"20",
		X"40",X"00",X"00",X"40",X"48",X"20",X"80",X"08",X"F8",X"08",X"88",X"40",X"88",X"08",X"60",X"60",
		X"20",X"78",X"20",X"20",X"B0",X"F8",X"48",X"80",X"48",X"80",X"80",X"88",X"88",X"20",X"08",X"A0",
		X"80",X"88",X"88",X"88",X"80",X"A8",X"A0",X"10",X"20",X"88",X"50",X"A8",X"50",X"20",X"40",X"40",
		X"10",X"08",X"00",X"00",X"FE",X"20",X"78",X"A8",X"88",X"F8",X"F0",X"BA",X"7C",X"20",X"44",X"44",
		X"6C",X"82",X"FF",X"FE",X"00",X"00",X"00",X"50",X"28",X"98",X"90",X"00",X"20",X"20",X"00",X"20",
		X"40",X"00",X"00",X"80",X"48",X"20",X"80",X"88",X"10",X"88",X"88",X"80",X"88",X"10",X"60",X"20",
		X"10",X"00",X"40",X"00",X"80",X"88",X"48",X"88",X"48",X"80",X"80",X"88",X"88",X"20",X"88",X"90",
		X"88",X"88",X"88",X"88",X"80",X"90",X"90",X"88",X"20",X"88",X"20",X"A8",X"88",X"20",X"80",X"40",
		X"08",X"08",X"00",X"00",X"48",X"20",X"F0",X"70",X"70",X"70",X"60",X"44",X"6C",X"50",X"38",X"82",
		X"00",X"82",X"FF",X"FE",X"00",X"20",X"00",X"50",X"F8",X"98",X"68",X"00",X"10",X"40",X"00",X"00",
		X"80",X"00",X"80",X"80",X"30",X"70",X"F8",X"70",X"10",X"70",X"70",X"80",X"70",X"60",X"00",X"40",
		X"00",X"00",X"00",X"20",X"78",X"88",X"F0",X"70",X"F0",X"F8",X"80",X"78",X"88",X"70",X"70",X"88",
		X"F8",X"88",X"88",X"F8",X"80",X"68",X"88",X"70",X"20",X"70",X"20",X"50",X"88",X"20",X"F8",X"70",
		X"08",X"70",X"00",X"F8",X"00",X"20",X"60",X"20",X"00",X"00",X"00",X"38",X"82",X"88",X"00",X"00",
		X"00",X"FE",X"FF",X"FE",X"00",X"11",X"41",X"30",X"21",X"10",X"20",X"31",X"00",X"01",X"03",X"06",
		X"0A",X"0F",X"15",X"1C",X"24",X"2D",X"08",X"10",X"08",X"10",X"0B",X"08",X"10",X"0D",X"0A",X"08",
		X"10",X"0E",X"0B",X"09",X"08",X"10",X"0E",X"0C",X"0A",X"09",X"08",X"10",X"0E",X"0D",X"0B",X"0A",
		X"09",X"08",X"10",X"0F",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"10",X"0F",X"0E",X"0C",X"0B",X"0A",
		X"09",X"09",X"08",X"10",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"09",X"08",X"00",X"19",X"32",
		X"4A",X"62",X"79",X"8E",X"A2",X"B5",X"C6",X"D5",X"E2",X"ED",X"F5",X"FB",X"FF",X"FF",X"FF",X"FB",
		X"F5",X"ED",X"E2",X"D5",X"C6",X"B5",X"A2",X"8E",X"79",X"62",X"4A",X"32",X"19",X"03",X"BD",X"03",
		X"87",X"03",X"54",X"03",X"24",X"02",X"F7",X"02",X"CD",X"02",X"A4",X"02",X"7E",X"02",X"5B",X"02",
		X"39",X"02",X"19",X"01",X"FB",X"01",X"DE",X"01",X"C3",X"01",X"AA",X"01",X"92",X"01",X"7C",X"01",
		X"66",X"01",X"52",X"01",X"3F",X"01",X"2D",X"01",X"1C",X"01",X"0C",X"00",X"FD",X"00",X"EF",X"00",
		X"E2",X"00",X"D5",X"00",X"C9",X"00",X"BE",X"00",X"B3",X"00",X"A9",X"00",X"A0",X"00",X"97",X"00",
		X"8E",X"00",X"86",X"00",X"7F",X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",
		X"5A",X"00",X"55",X"00",X"50",X"00",X"4B",X"00",X"47",X"00",X"43",X"00",X"3F",X"00",X"3C",X"00",
		X"38",X"00",X"35",X"00",X"32",X"00",X"2F",X"00",X"2D",X"00",X"2A",X"00",X"28",X"00",X"26",X"00",
		X"24",X"00",X"22",X"00",X"20",X"00",X"1E",X"00",X"1C",X"00",X"1B",X"00",X"00",X"FE",X"E8",X"FE",
		X"B6",X"93",X"1F",X"0C",X"93",X"1F",X"06",X"98",X"9F",X"24",X"3C",X"11",X"80",X"FD",X"69",X"FD",
		X"79",X"21",X"07",X"21",X"07",X"21",X"07",X"21",X"07",X"21",X"07",X"21",X"07",X"21",X"0E",X"99",
		X"9F",X"24",X"0E",X"95",X"9B",X"20",X"0E",X"21",X"07",X"21",X"07",X"21",X"07",X"21",X"07",X"21",
		X"07",X"21",X"07",X"9D",X"A3",X"28",X"0E",X"A0",X"A6",X"2B",X"0E",X"22",X"02",X"28",X"02",X"2D",
		X"02",X"28",X"02",X"22",X"02",X"28",X"02",X"2D",X"02",X"28",X"02",X"22",X"02",X"28",X"02",X"2D",
		X"02",X"28",X"02",X"2E",X"02",X"2D",X"28",X"21",X"80",X"EF",X"FF",X"FE",X"DC",X"BA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"01",X"00",X"FF",X"FE",
		X"FF",X"FD",X"C3",X"FE",X"B6",X"51",X"24",X"50",X"06",X"50",X"06",X"50",X"0C",X"50",X"06",X"50",
		X"06",X"50",X"04",X"50",X"04",X"50",X"04",X"50",X"18",X"50",X"04",X"50",X"04",X"50",X"04",X"50",
		X"0C",X"50",X"0C",X"50",X"24",X"50",X"06",X"50",X"06",X"50",X"0C",X"50",X"06",X"50",X"06",X"50",
		X"04",X"50",X"04",X"50",X"04",X"50",X"18",X"50",X"04",X"50",X"04",X"50",X"04",X"50",X"0C",X"50",
		X"18",X"26",X"80",X"FD",X"BA",X"98",X"76",X"55",X"44",X"33",X"22",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FE",X"28",X"FD",X"79",X"98",X"1C",X"10",X"3F",X"08",X"98",X"1C",X"04",X"98",
		X"1C",X"04",X"98",X"1C",X"10",X"3F",X"08",X"98",X"1C",X"04",X"98",X"1C",X"04",X"98",X"1C",X"08",
		X"93",X"18",X"08",X"98",X"1C",X"08",X"9C",X"1F",X"08",X"98",X"1C",X"08",X"93",X"18",X"08",X"98",
		X"1C",X"08",X"93",X"18",X"08",X"98",X"1C",X"08",X"9C",X"1F",X"08",X"98",X"1C",X"08",X"93",X"18",
		X"08",X"98",X"1C",X"08",X"93",X"18",X"08",X"98",X"1C",X"08",X"9C",X"1F",X"08",X"98",X"1C",X"08",
		X"93",X"18",X"08",X"9C",X"1F",X"30",X"1A",X"80",X"FF",X"FE",X"DC",X"BA",X"98",X"76",X"54",X"32",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"66",X"FE",X"B6",X"0C",X"18",X"11",X"18",
		X"0C",X"18",X"11",X"18",X"0C",X"18",X"11",X"18",X"0C",X"12",X"0C",X"06",X"11",X"18",X"9D",X"21",
		X"18",X"9F",X"23",X"18",X"A1",X"24",X"18",X"A3",X"26",X"18",X"9F",X"A4",X"28",X"18",X"07",X"12",
		X"07",X"06",X"00",X"3C",X"18",X"80",X"DE",X"EF",X"FE",X"DC",X"BA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"B2",X"FE",X"B6",X"18",X"06",X"1A",X"06",X"1C",X"0C",
		X"18",X"0C",X"1A",X"24",X"23",X"18",X"17",X"06",X"18",X"06",X"1A",X"0C",X"17",X"0C",X"18",X"24",
		X"24",X"18",X"A4",X"28",X"0C",X"A3",X"26",X"0C",X"A1",X"24",X"0C",X"9F",X"23",X"0C",X"9D",X"21",
		X"18",X"9A",X"1F",X"18",X"17",X"06",X"18",X"06",X"1A",X"0C",X"17",X"0C",X"18",X"24",X"24",X"24",
		X"18",X"80",X"FF",X"EE",X"DD",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"E8",X"FE",X"B6",X"96",X"9A",X"1D",X"1E",X"91",X"95",
		X"18",X"1E",X"94",X"98",X"1B",X"1E",X"8F",X"94",X"18",X"14",X"16",X"0A",X"8C",X"91",X"15",X"14",
		X"16",X"0A",X"91",X"95",X"18",X"32",X"18",X"80",X"EE",X"FF",X"FF",X"EE",X"EE",X"DD",X"CC",X"BB",
		X"AA",X"99",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"16",X"FE",X"B6",X"1C",X"06",X"1F",X"06",
		X"1C",X"06",X"18",X"06",X"1A",X"06",X"18",X"06",X"15",X"06",X"13",X"06",X"18",X"06",X"13",X"06",
		X"17",X"06",X"18",X"1E",X"18",X"80",X"FF",X"FF",X"EE",X"EE",X"DD",X"DD",X"CC",X"CC",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"28",X"FE",X"B6",X"16",X"0F",X"16",X"05",X"16",X"05",
		X"16",X"05",X"1A",X"0F",X"16",X"0F",X"1D",X"0F",X"1D",X"05",X"1D",X"05",X"1D",X"05",X"21",X"0F",
		X"1D",X"32",X"1D",X"80",X"FE",X"28",X"FE",X"B6",X"16",X"06",X"16",X"02",X"16",X"02",X"16",X"02",
		X"1A",X"06",X"16",X"06",X"1D",X"06",X"1D",X"02",X"1D",X"02",X"1D",X"02",X"21",X"06",X"1D",X"32",
		X"11",X"80",X"FE",X"28",X"FE",X"B6",X"1B",X"0F",X"16",X"05",X"16",X"05",X"16",X"05",X"17",X"30",
		X"16",X"05",X"16",X"05",X"16",X"05",X"17",X"30",X"16",X"80",X"FD",X"69",X"FE",X"B6",X"A0",X"23",
		X"12",X"A0",X"23",X"0C",X"9C",X"20",X"06",X"9E",X"21",X"12",X"9C",X"20",X"32",X"13",X"80",X"FD",
		X"C3",X"FE",X"B6",X"16",X"04",X"16",X"04",X"16",X"04",X"16",X"04",X"1A",X"08",X"1C",X"80",X"A6",
		X"A0",X"20",X"08",X"BD",X"F3",X"BE",X"B6",X"C8",X"80",X"84",X"7F",X"B7",X"C8",X"80",X"7A",X"C8",
		X"80",X"A6",X"A4",X"47",X"84",X"F8",X"E6",X"A0",X"58",X"58",X"58",X"58",X"57",X"C4",X"F8",X"7D",
		X"C8",X"80",X"2B",X"DF",X"BD",X"F3",X"DF",X"B6",X"C8",X"80",X"85",X"0F",X"26",X"E0",X"85",X"20",
		X"27",X"CD",X"39",X"4B",X"41",X"52",X"52",X"53",X"4F",X"46",X"54",X"38",X"32",X"4C",X"44",X"4D",
		X"43",X"42",X"43",X"4A",X"54",X"38",X"32",X"4C",X"44",X"4D",X"43",X"42",X"43",X"4A",X"00",X"00",
		X"00",X"00",X"CB",X"F2",X"CB",X"F2",X"CB",X"F5",X"CB",X"F8",X"CB",X"FB",X"CB",X"FB",X"F0",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
