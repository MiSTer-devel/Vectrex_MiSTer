--------------------------------------------------------------------------------
-- VECTREX
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- DO 8/2017
--------------------------------------------------------------------------------

-- EXECUTIVE ROM

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

USE std.textio.ALL;

LIBRARY work;
USE work.base_pack.ALL;
USE work.mc6809_pack.ALL;
USE work.plomb_pack.ALL;
USE work.vid_pack.ALL;

ENTITY exerom IS
  PORT (
    ad  : IN uv16;
    dr  : OUT uv8;
    clk : IN std_logic
    );
END ENTITY exerom;


ARCHITECTURE rtl OF exerom IS

  -- EXECUTIVE
  CONSTANT rom: arr_uv8 := (
    x"ed",x"77",x"f8",x"50",x"30",x"e8",x"4d",x"49",x"4e",x"45",x"80",x"f8",
    x"50",x"00",x"de",x"53",x"54",x"4f",x"52",x"4d",x"80",x"00",x"8e",x"c8",
    x"83",x"6f",x"80",x"8c",x"cb",x"c5",x"26",x"f9",x"bd",x"e8",x"e3",x"7c",
    x"c8",x"24",x"86",x"bb",x"b7",x"c8",x"80",x"8e",x"01",x"01",x"bf",x"c8",
    x"81",x"8e",x"c8",x"83",x"6f",x"80",x"8c",x"cb",x"70",x"26",x"f9",x"20",
    x"00",x"bd",x"f1",x"af",x"cc",x"02",x"00",x"bd",x"f7",x"a9",x"0a",x"79",
    x"0f",x"56",x"0f",x"9b",x"8e",x"c8",x"a8",x"bd",x"f8",x"4f",x"8e",x"c8",
    x"af",x"bd",x"f8",x"4f",x"8e",x"c8",x"f9",x"bd",x"f8",x"4f",x"cc",x"00",
    x"01",x"bd",x"f8",x"7c",x"8e",x"c9",x"00",x"bd",x"f8",x"4f",x"cc",x"00",
    x"01",x"bd",x"f8",x"7c",x"8e",x"ed",x"ab",x"9f",x"c4",x"9f",x"c6",x"86",
    x"05",x"97",x"d9",x"97",x"da",x"97",x"db",x"20",x"24",x"bd",x"e8",x"66",
    x"10",x"8e",x"c8",x"c4",x"96",x"9b",x"ae",x"a6",x"30",x"04",x"af",x"a6",
    x"8e",x"ed",x"a7",x"96",x"9b",x"ae",x"86",x"a6",x"05",x"84",x"03",x"26",
    x"02",x"0c",x"d9",x"cc",x"00",x"01",x"bd",x"f8",x"7c",x"bd",x"e7",x"e4",
    x"8e",x"c8",x"c4",x"96",x"9b",x"ae",x"86",x"a6",x"84",x"2b",x"05",x"bd",
    x"e1",x"29",x"20",x"41",x"dc",x"f0",x"83",x"00",x"01",x"dd",x"f0",x"27",
    x"14",x"34",x"08",x"bd",x"f1",x"aa",x"bd",x"ea",x"cf",x"ce",x"ee",x"2f",
    x"bd",x"ea",x"9d",x"35",x"08",x"96",x"0f",x"27",x"24",x"8e",x"c8",x"a8",
    x"ce",x"cb",x"eb",x"bd",x"f8",x"d8",x"8e",x"c8",x"af",x"ce",x"cb",x"eb",
    x"bd",x"f8",x"d8",x"dc",x"f0",x"10",x"26",x"ff",x"44",x"bd",x"f1",x"8b",
    x"0f",x"3b",x"10",x"ce",x"cb",x"ea",x"7e",x"f0",x"1c",x"34",x"08",x"bd",
    x"ea",x"f0",x"bd",x"e5",x"1e",x"bd",x"e2",x"62",x"bd",x"e4",x"b8",x"bd",
    x"e3",x"53",x"35",x"08",x"bd",x"eb",x"43",x"bd",x"ec",x"46",x"bd",x"ec",
    x"95",x"bd",x"e6",x"47",x"25",x"df",x"96",x"bd",x"10",x"27",x"ff",x"61",
    x"96",x"be",x"10",x"26",x"ff",x"92",x"7e",x"e0",x"a5",x"9f",x"c2",x"cc",
    x"7f",x"00",x"dd",x"dc",x"97",x"b7",x"86",x"20",x"97",x"9c",x"8e",x"e1",
    x"e7",x"9f",x"9d",x"8e",x"c9",x"33",x"9f",x"b9",x"86",x"1d",x"97",x"b8",
    x"0f",x"56",x"ce",x"ed",x"77",x"bd",x"f6",x"8d",x"34",x"08",x"bd",x"e7",
    x"11",x"bd",x"f6",x"87",x"96",x"26",x"85",x"01",x"26",x"02",x"0a",x"b7",
    x"bd",x"ea",x"f0",x"bd",x"ea",x"cf",x"bd",x"f2",x"89",x"bd",x"e5",x"1e",
    x"bd",x"f2",x"a5",x"f6",x"c8",x"b7",x"27",x"1c",x"8e",x"ef",x"26",x"10",
    x"be",x"c8",x"dc",x"bd",x"ea",x"7f",x"8e",x"ef",x"5d",x"bd",x"ea",x"7f",
    x"8e",x"ef",x"94",x"bd",x"ea",x"7f",x"35",x"08",x"0a",x"dc",x"20",x"c0",
    x"35",x"08",x"0f",x"9c",x"86",x"04",x"97",x"b7",x"86",x"7f",x"97",x"b8",
    x"96",x"b7",x"27",x"4a",x"d6",x"b8",x"27",x"04",x"0a",x"b8",x"20",x"12",
    x"d6",x"26",x"c4",x"1f",x"26",x"0c",x"4a",x"97",x"b7",x"9e",x"c2",x"a6",
    x"86",x"c6",x"03",x"bd",x"e9",x"a1",x"34",x"08",x"bd",x"ea",x"f0",x"bd",
    x"f2",x"a9",x"ce",x"ee",x"20",x"bd",x"ea",x"9d",x"10",x"8e",x"e0",x"f8",
    x"ce",x"ed",x"a7",x"b6",x"c8",x"9b",x"ee",x"c6",x"bd",x"ea",x"a8",x"bd",
    x"e5",x"1e",x"bd",x"e2",x"62",x"bd",x"e4",x"b8",x"35",x"08",x"bd",x"eb",
    x"43",x"bd",x"e6",x"47",x"20",x"b2",x"39",x"0a",x"b8",x"27",x"4e",x"0c",
    x"ed",x"bd",x"f5",x"17",x"84",x"07",x"8b",x"04",x"97",x"9c",x"de",x"b9",
    x"86",x"80",x"a7",x"c4",x"dc",x"dc",x"8b",x"08",x"a7",x"44",x"6f",x"45",
    x"e7",x"46",x"6f",x"47",x"bd",x"f5",x"17",x"4d",x"2b",x"0c",x"81",x"10",
    x"2c",x"02",x"8b",x"0c",x"81",x"60",x"2f",x"0e",x"20",x"ee",x"81",x"f0",
    x"2f",x"02",x"80",x"0c",x"81",x"a0",x"2c",x"02",x"20",x"e2",x"a7",x"c8",
    x"11",x"1f",x"89",x"1d",x"8a",x"01",x"a7",x"c8",x"10",x"6f",x"42",x"31",
    x"c8",x"12",x"10",x"9f",x"b9",x"39",x"00",x"02",x"07",x"10",x"00",x"20",
    x"18",x"10",x"01",x"00",x"05",x"00",x"03",x"25",x"07",x"50",x"00",x"00",
    x"01",x"00",x"00",x"35",x"00",x"00",x"00",x"00",x"04",x"04",x"08",x"08",
    x"0d",x"0d",x"ee",x"3d",x"ee",x"53",x"ee",x"6f",x"ee",x"8e",x"34",x"08",
    x"86",x"c8",x"1f",x"8b",x"96",x"bd",x"10",x"26",x"00",x"9c",x"96",x"ee",
    x"10",x"26",x"00",x"a7",x"96",x"13",x"10",x"26",x"00",x"92",x"96",x"14",
    x"27",x"32",x"96",x"d4",x"91",x"d6",x"27",x"1c",x"91",x"d8",x"27",x"08",
    x"96",x"d5",x"27",x"14",x"96",x"d7",x"26",x"20",x"96",x"d7",x"8b",x"0c",
    x"81",x"7f",x"22",x"18",x"97",x"d7",x"96",x"d4",x"97",x"d8",x"20",x"0e",
    x"96",x"d5",x"8b",x"0c",x"81",x"7f",x"22",x"08",x"97",x"d5",x"96",x"d4",
    x"97",x"d6",x"0c",x"f2",x"96",x"d5",x"27",x"0e",x"80",x"02",x"97",x"d5",
    x"d6",x"d6",x"bd",x"e7",x"b5",x"10",x"9f",x"cc",x"9f",x"ce",x"96",x"d7",
    x"27",x"0e",x"80",x"02",x"97",x"d7",x"d6",x"d8",x"bd",x"e7",x"b5",x"10",
    x"9f",x"d0",x"9f",x"d2",x"dc",x"c8",x"d3",x"cc",x"d3",x"d0",x"dd",x"c8",
    x"dc",x"ca",x"d3",x"ce",x"d3",x"d2",x"dd",x"ca",x"96",x"1b",x"27",x"0f",
    x"2b",x"04",x"0a",x"d4",x"20",x"06",x"0c",x"d4",x"20",x"02",x"34",x"08",
    x"bd",x"e8",x"4c",x"86",x"d0",x"1f",x"8b",x"bd",x"f2",x"a5",x"c6",x"0c",
    x"10",x"8e",x"c8",x"c8",x"8e",x"cb",x"89",x"bd",x"ea",x"8d",x"35",x"88",
    x"86",x"80",x"97",x"ee",x"bd",x"f5",x"17",x"84",x"03",x"8b",x"03",x"97",
    x"ef",x"0c",x"f6",x"96",x"ee",x"2a",x"19",x"0a",x"ef",x"27",x"0d",x"bd",
    x"e9",x"8a",x"97",x"c8",x"0f",x"c9",x"d7",x"ca",x"0f",x"cb",x"35",x"88",
    x"04",x"ee",x"86",x"1f",x"97",x"ef",x"35",x"88",x"d6",x"ef",x"c1",x"e0",
    x"2f",x"0c",x"96",x"ef",x"80",x"04",x"97",x"ef",x"4f",x"bd",x"e9",x"4a",
    x"35",x"88",x"0f",x"ef",x"0f",x"ee",x"bd",x"e8",x"37",x"35",x"88",x"b6",
    x"c8",x"e7",x"27",x"2b",x"34",x"08",x"86",x"c8",x"1f",x"8b",x"96",x"e7",
    x"27",x"21",x"dc",x"de",x"d3",x"e2",x"dd",x"de",x"97",x"dc",x"dc",x"e0",
    x"d3",x"e4",x"dd",x"e0",x"97",x"dd",x"35",x"08",x"bd",x"f2",x"a5",x"c6",
    x"08",x"10",x"be",x"c8",x"dc",x"8e",x"ef",x"b3",x"bd",x"ea",x"7f",x"39",
    x"8e",x"e3",x"a1",x"9f",x"a3",x"bd",x"f5",x"17",x"8e",x"e4",x"48",x"84",
    x"06",x"ae",x"86",x"ec",x"81",x"dd",x"dc",x"97",x"de",x"0f",x"df",x"d7",
    x"e0",x"0f",x"e1",x"20",x"58",x"96",x"bf",x"26",x"19",x"bd",x"f5",x"17",
    x"84",x"7f",x"8b",x"30",x"97",x"a2",x"bd",x"f5",x"17",x"84",x"3f",x"97",
    x"e6",x"bd",x"f5",x"17",x"8b",x"10",x"97",x"e7",x"20",x"49",x"96",x"bd",
    x"26",x"e3",x"c6",x"1c",x"ce",x"c9",x"33",x"a6",x"c4",x"27",x"08",x"33",
    x"c8",x"12",x"5a",x"26",x"f6",x"20",x"34",x"0c",x"ed",x"0a",x"bf",x"9e",
    x"de",x"af",x"44",x"9e",x"e0",x"af",x"46",x"86",x"40",x"a7",x"c4",x"96",
    x"c0",x"26",x"10",x"8e",x"e4",x"12",x"9f",x"9d",x"bd",x"f5",x"17",x"84",
    x"7f",x"8b",x"40",x"97",x"9c",x"0c",x"c0",x"9e",x"e8",x"a6",x"80",x"97",
    x"a2",x"a6",x"80",x"97",x"e6",x"a6",x"80",x"97",x"e7",x"9f",x"e8",x"d6",
    x"e6",x"bd",x"e7",x"b5",x"10",x"9f",x"e2",x"9f",x"e4",x"39",x"ce",x"c8",
    x"c4",x"96",x"9b",x"ee",x"c6",x"a6",x"c4",x"c6",x"03",x"bd",x"e9",x"a1",
    x"8e",x"e4",x"26",x"9f",x"9d",x"39",x"0a",x"c1",x"27",x"06",x"86",x"ff",
    x"97",x"9c",x"20",x"17",x"bd",x"f5",x"17",x"1f",x"89",x"c4",x"03",x"26",
    x"02",x"cb",x"01",x"ce",x"c8",x"c4",x"96",x"9b",x"ee",x"c6",x"a6",x"c4",
    x"bd",x"e9",x"a1",x"39",x"e4",x"50",x"e4",x"6a",x"e4",x"84",x"e4",x"9e",
    x"7f",x"00",x"28",x"20",x"30",x"40",x"28",x"30",x"28",x"00",x"10",x"30",
    x"10",x"40",x"18",x"20",x"50",x"40",x"30",x"28",x"30",x"08",x"60",x"7f",
    x"38",x"70",x"80",x"00",x"40",x"00",x"30",x"20",x"10",x"50",x"20",x"28",
    x"40",x"30",x"3e",x"70",x"18",x"30",x"60",x"20",x"18",x"40",x"30",x"24",
    x"50",x"7f",x"06",x"70",x"00",x"7f",x"40",x"10",x"60",x"28",x"38",x"30",
    x"28",x"08",x"40",x"30",x"28",x"7f",x"20",x"18",x"30",x"30",x"08",x"68",
    x"40",x"20",x"50",x"7f",x"38",x"70",x"00",x"80",x"40",x"30",x"60",x"38",
    x"18",x"30",x"30",x"20",x"18",x"20",x"38",x"40",x"28",x"10",x"60",x"20",
    x"00",x"30",x"40",x"38",x"50",x"7f",x"1c",x"70",x"86",x"04",x"ce",x"c9",
    x"0b",x"8e",x"c8",x"15",x"b7",x"c8",x"8f",x"bd",x"f2",x"a9",x"a6",x"c4",
    x"27",x"22",x"6a",x"49",x"27",x"19",x"ec",x"45",x"e3",x"41",x"ed",x"45",
    x"ec",x"47",x"e3",x"43",x"ed",x"47",x"31",x"45",x"bd",x"ea",x"6d",x"33",
    x"4a",x"7a",x"c8",x"8f",x"26",x"e0",x"39",x"6f",x"c4",x"7a",x"c8",x"ea",
    x"b6",x"c8",x"bd",x"26",x"ee",x"b6",x"c8",x"ee",x"26",x"e9",x"a6",x"84",
    x"27",x"e5",x"6f",x"84",x"7c",x"c8",x"b6",x"6c",x"c4",x"fc",x"c8",x"c8",
    x"ed",x"45",x"fc",x"c8",x"ca",x"ed",x"47",x"fc",x"c9",x"07",x"ed",x"41",
    x"fc",x"c9",x"09",x"ed",x"43",x"86",x"18",x"a7",x"49",x"7c",x"c8",x"ea",
    x"20",x"c1",x"86",x"1c",x"b7",x"c8",x"8f",x"ce",x"c9",x"33",x"a6",x"c4",
    x"26",x"09",x"33",x"c8",x"12",x"7a",x"c8",x"8f",x"26",x"f4",x"39",x"10",
    x"2b",x"00",x"9c",x"85",x"40",x"10",x"26",x"00",x"a4",x"85",x"20",x"10",
    x"26",x"00",x"a9",x"85",x"10",x"10",x"26",x"00",x"d4",x"85",x"01",x"10",
    x"26",x"00",x"d8",x"a6",x"41",x"81",x"04",x"27",x"56",x"85",x"01",x"27",
    x"31",x"b6",x"c8",x"ee",x"26",x"2c",x"b6",x"c8",x"bd",x"26",x"27",x"34",
    x"08",x"bd",x"f1",x"af",x"96",x"c8",x"a0",x"44",x"d6",x"ca",x"e0",x"46",
    x"bd",x"f5",x"93",x"80",x"10",x"97",x"83",x"8e",x"e2",x"3e",x"e6",x"43",
    x"a6",x"85",x"d6",x"83",x"bd",x"e7",x"b5",x"10",x"af",x"48",x"af",x"4a",
    x"35",x"08",x"ec",x"44",x"e3",x"48",x"ed",x"44",x"ec",x"46",x"e3",x"4a",
    x"ed",x"46",x"bd",x"f2",x"a5",x"8e",x"e2",x"5a",x"a6",x"41",x"48",x"ae",
    x"86",x"31",x"44",x"e6",x"42",x"bd",x"ea",x"8d",x"7e",x"e5",x"2a",x"ec",
    x"44",x"e3",x"48",x"29",x"1a",x"ed",x"44",x"ec",x"46",x"e3",x"4a",x"29",
    x"12",x"ed",x"46",x"bd",x"f2",x"a9",x"31",x"44",x"8e",x"cb",x"a7",x"c6",
    x"04",x"bd",x"ea",x"8d",x"7e",x"e5",x"2a",x"6f",x"c4",x"7a",x"c8",x"eb",
    x"7e",x"e5",x"2a",x"a6",x"46",x"ab",x"c8",x"10",x"a7",x"46",x"a1",x"c8",
    x"11",x"26",x"02",x"64",x"c4",x"bd",x"f2",x"a5",x"31",x"44",x"bd",x"ea",
    x"6d",x"7e",x"e5",x"2a",x"a6",x"43",x"81",x"03",x"26",x"0d",x"a6",x"42",
    x"a1",x"c8",x"10",x"2c",x"06",x"8b",x"08",x"a7",x"42",x"20",x"1b",x"64",
    x"c4",x"a6",x"c8",x"10",x"a7",x"42",x"86",x"18",x"a7",x"c8",x"10",x"b6",
    x"c8",x"ed",x"26",x"0a",x"b6",x"c8",x"c0",x"26",x"05",x"86",x"7f",x"b7",
    x"c8",x"a2",x"7e",x"e5",x"96",x"6a",x"c8",x"10",x"26",x"02",x"64",x"c4",
    x"7e",x"e5",x"96",x"6f",x"c4",x"a6",x"41",x"81",x"04",x"27",x"15",x"e6",
    x"43",x"5a",x"27",x"10",x"34",x"0a",x"86",x"c8",x"1f",x"8b",x"a6",x"e4",
    x"bd",x"e9",x"a1",x"bd",x"e9",x"a1",x"35",x"0a",x"7e",x"e5",x"2a",x"34",
    x"08",x"bd",x"f1",x"aa",x"bd",x"f2",x"a9",x"ce",x"cb",x"2b",x"86",x"0e",
    x"b7",x"c8",x"8f",x"a6",x"c4",x"10",x"27",x"00",x"a6",x"e6",x"44",x"e1",
    x"41",x"24",x"0d",x"cb",x"03",x"e7",x"44",x"10",x"ae",x"42",x"8e",x"ee",
    x"ba",x"bd",x"ea",x"7f",x"4d",x"10",x"2a",x"00",x"83",x"7a",x"c8",x"f7",
    x"10",x"27",x"00",x"37",x"b6",x"c8",x"26",x"84",x"01",x"26",x"03",x"7c",
    x"c8",x"f8",x"b6",x"c8",x"f8",x"10",x"8e",x"7f",x"00",x"8e",x"ef",x"04",
    x"bd",x"e7",x"6a",x"10",x"8e",x"60",x"80",x"8e",x"ef",x"0b",x"bd",x"e7",
    x"6a",x"10",x"8e",x"80",x"50",x"8e",x"ef",x"15",x"bd",x"e7",x"6a",x"10",
    x"8e",x"a0",x"80",x"8e",x"ef",x"1c",x"bd",x"e7",x"6a",x"20",x"50",x"7a",
    x"c8",x"d9",x"7f",x"c8",x"eb",x"7f",x"c8",x"ed",x"b6",x"c8",x"79",x"27",
    x"2b",x"b6",x"c8",x"9b",x"44",x"8e",x"c8",x"da",x"f6",x"c8",x"d9",x"e7",
    x"86",x"b6",x"c8",x"da",x"26",x"05",x"b6",x"c8",x"db",x"27",x"1a",x"b6",
    x"c8",x"9b",x"8b",x"02",x"84",x"02",x"b7",x"c8",x"9b",x"44",x"8e",x"c8",
    x"da",x"e6",x"86",x"f7",x"c8",x"d9",x"27",x"eb",x"b6",x"c8",x"d9",x"26",
    x"0d",x"86",x"01",x"b7",x"c8",x"be",x"20",x"06",x"e6",x"44",x"e1",x"41",
    x"25",x"05",x"6f",x"c4",x"7a",x"c8",x"ec",x"33",x"45",x"7a",x"c8",x"8f",
    x"10",x"26",x"ff",x"4b",x"bd",x"ec",x"c9",x"20",x"05",x"34",x"08",x"bd",
    x"f1",x"aa",x"bd",x"f2",x"a5",x"8e",x"80",x"38",x"bf",x"c8",x"90",x"b6",
    x"c8",x"d9",x"27",x"1e",x"b7",x"c8",x"8f",x"7a",x"c8",x"8f",x"27",x"16",
    x"b6",x"c8",x"91",x"8b",x"06",x"b7",x"c8",x"91",x"c6",x"04",x"10",x"be",
    x"c8",x"90",x"8e",x"ee",x"eb",x"bd",x"ea",x"7f",x"20",x"e5",x"35",x"08",
    x"96",x"26",x"84",x"01",x"48",x"48",x"48",x"8e",x"ee",x"ad",x"ce",x"cb",
    x"a7",x"bd",x"f6",x"1f",x"d6",x"ec",x"26",x"0f",x"96",x"bd",x"26",x"08",
    x"d6",x"eb",x"26",x"07",x"d6",x"ed",x"26",x"03",x"1c",x"fe",x"39",x"1a",
    x"01",x"39",x"34",x"32",x"8e",x"c8",x"c8",x"bd",x"f2",x"f2",x"a6",x"e4",
    x"97",x"04",x"1f",x"20",x"bd",x"f3",x"12",x"c6",x"0c",x"ae",x"61",x"bd",
    x"f4",x"0e",x"35",x"b2",x"34",x"16",x"8e",x"cb",x"2b",x"86",x"0e",x"e6",
    x"84",x"27",x"07",x"30",x"05",x"4a",x"26",x"f7",x"20",x"1d",x"a6",x"e4",
    x"84",x"80",x"4c",x"a7",x"84",x"2a",x"02",x"0c",x"bd",x"a6",x"e4",x"84",
    x"7f",x"a7",x"04",x"a6",x"61",x"a7",x"01",x"ec",x"62",x"ed",x"02",x"0c",
    x"ec",x"0c",x"f3",x"35",x"96",x"34",x"36",x"bd",x"f6",x"01",x"a7",x"64",
    x"1d",x"58",x"49",x"58",x"49",x"58",x"49",x"ed",x"62",x"e6",x"64",x"1d",
    x"58",x"49",x"58",x"49",x"58",x"49",x"ed",x"64",x"35",x"b6",x"34",x"36",
    x"8d",x"df",x"ec",x"7c",x"58",x"49",x"ed",x"64",x"ec",x"7a",x"58",x"49",
    x"ed",x"62",x"35",x"b6",x"86",x"d0",x"1f",x"8b",x"bd",x"f2",x"72",x"86",
    x"c8",x"1f",x"8b",x"0f",x"9c",x"0f",x"9f",x"0f",x"a2",x"0f",x"a5",x"8e",
    x"c9",x"0b",x"6f",x"80",x"8c",x"cb",x"71",x"26",x"f9",x"cc",x"00",x"00",
    x"dd",x"de",x"dd",x"e0",x"dd",x"e2",x"dd",x"e4",x"97",x"e7",x"97",x"bd",
    x"97",x"be",x"97",x"ea",x"97",x"eb",x"97",x"ec",x"97",x"f8",x"c6",x"40",
    x"d7",x"f7",x"97",x"ed",x"97",x"c0",x"8e",x"08",x"00",x"9f",x"f0",x"86",
    x"07",x"97",x"bf",x"8e",x"e3",x"84",x"9f",x"a3",x"cc",x"00",x"00",x"dd",
    x"c8",x"dd",x"ca",x"cc",x"00",x"00",x"97",x"d4",x"dd",x"cc",x"dd",x"ce",
    x"97",x"d5",x"97",x"d6",x"dd",x"d0",x"dd",x"d2",x"97",x"d7",x"97",x"d8",
    x"96",x"d4",x"8e",x"ee",x"eb",x"ce",x"cb",x"89",x"bd",x"f6",x"1f",x"86",
    x"7f",x"d6",x"d4",x"bd",x"e7",x"d2",x"10",x"bf",x"c9",x"07",x"bf",x"c9",
    x"09",x"39",x"34",x"30",x"34",x"08",x"bd",x"f1",x"aa",x"bd",x"f2",x"72",
    x"35",x"08",x"86",x"a0",x"97",x"8f",x"96",x"c8",x"27",x"0a",x"2b",x"03",
    x"4a",x"20",x"01",x"4c",x"97",x"c8",x"0f",x"c9",x"96",x"ca",x"27",x"0a",
    x"2b",x"03",x"4a",x"20",x"01",x"4c",x"97",x"ca",x"0f",x"cb",x"96",x"d4",
    x"27",x"0c",x"81",x"1f",x"2e",x"03",x"4a",x"20",x"01",x"4c",x"84",x"3f",
    x"97",x"d4",x"bd",x"e2",x"f2",x"8e",x"cb",x"81",x"c6",x"08",x"a6",x"84",
    x"8b",x"03",x"a7",x"80",x"5a",x"26",x"f7",x"34",x"08",x"bd",x"f1",x"aa",
    x"bd",x"ea",x"cf",x"5f",x"86",x"20",x"bd",x"e9",x"0b",x"bd",x"e8",x"fd",
    x"35",x"08",x"96",x"c8",x"10",x"26",x"ff",x"aa",x"96",x"ca",x"10",x"26",
    x"ff",x"a4",x"96",x"d4",x"10",x"26",x"ff",x"9e",x"0a",x"8f",x"10",x"26",
    x"ff",x"98",x"bd",x"e7",x"e4",x"35",x"b0",x"8e",x"ed",x"e0",x"10",x"8e",
    x"cb",x"71",x"ce",x"cb",x"81",x"c6",x"08",x"86",x"16",x"af",x"a1",x"30",
    x"08",x"a7",x"c0",x"8b",x"0f",x"5a",x"26",x"f5",x"39",x"34",x"1e",x"8e",
    x"cb",x"81",x"86",x"08",x"6c",x"80",x"4a",x"26",x"fb",x"20",x"02",x"34",
    x"1e",x"86",x"d0",x"1f",x"8b",x"86",x"09",x"34",x"02",x"6a",x"e4",x"26",
    x"07",x"bd",x"f3",x"54",x"35",x"02",x"35",x"9e",x"bd",x"f3",x"54",x"86",
    x"03",x"b7",x"c8",x"23",x"a6",x"e4",x"4a",x"8e",x"cb",x"81",x"e6",x"86",
    x"c4",x"7f",x"e1",x"61",x"23",x"df",x"e0",x"62",x"2f",x"db",x"d7",x"04",
    x"8e",x"cb",x"71",x"48",x"ae",x"86",x"bd",x"f2",x"a9",x"bd",x"f2",x"d5",
    x"20",x"cb",x"34",x"1e",x"86",x"d0",x"1f",x"8b",x"86",x"09",x"34",x"02",
    x"6a",x"e4",x"26",x"07",x"bd",x"f3",x"54",x"35",x"02",x"35",x"9e",x"bd",
    x"f3",x"54",x"86",x"03",x"b7",x"c8",x"23",x"8e",x"c8",x"c8",x"bd",x"f2",
    x"f2",x"e6",x"e4",x"58",x"58",x"eb",x"62",x"2f",x"df",x"c4",x"7f",x"d7",
    x"04",x"8e",x"cb",x"71",x"a6",x"e4",x"4a",x"48",x"ae",x"86",x"bd",x"f2",
    x"a9",x"bd",x"f2",x"d5",x"20",x"ca",x"34",x"06",x"bd",x"f5",x"17",x"a7",
    x"e4",x"bd",x"f5",x"17",x"81",x"60",x"2e",x"f9",x"81",x"a0",x"2d",x"f5",
    x"a7",x"61",x"35",x"06",x"39",x"34",x"76",x"96",x"ed",x"10",x"27",x"00",
    x"93",x"0a",x"ed",x"bd",x"f5",x"17",x"84",x"1f",x"97",x"8b",x"81",x"1b",
    x"23",x"04",x"80",x"04",x"20",x"f6",x"c6",x"12",x"3d",x"c3",x"c9",x"33",
    x"1f",x"03",x"a6",x"c4",x"84",x"c0",x"26",x"0d",x"0c",x"8b",x"96",x"8b",
    x"81",x"1b",x"2f",x"ea",x"0f",x"8b",x"4f",x"20",x"e5",x"a6",x"e4",x"a7",
    x"41",x"8e",x"e2",x"42",x"48",x"10",x"ae",x"86",x"10",x"9f",x"89",x"c6",
    x"20",x"e7",x"c4",x"8e",x"e2",x"3e",x"a6",x"61",x"e6",x"86",x"d7",x"8b",
    x"8e",x"e2",x"3a",x"e6",x"86",x"e7",x"c8",x"10",x"a7",x"43",x"8e",x"e2",
    x"52",x"48",x"10",x"ae",x"86",x"10",x"af",x"4c",x"8e",x"e2",x"4a",x"10",
    x"ae",x"86",x"10",x"9f",x"87",x"81",x"06",x"26",x"02",x"0c",x"f4",x"96",
    x"88",x"9b",x"8a",x"19",x"a7",x"4f",x"96",x"87",x"99",x"89",x"19",x"a7",
    x"4e",x"96",x"8b",x"bd",x"ea",x"3e",x"bd",x"e7",x"b5",x"10",x"af",x"48",
    x"af",x"4a",x"0c",x"eb",x"96",x"c0",x"27",x"08",x"86",x"ff",x"97",x"9c",
    x"86",x"03",x"97",x"c1",x"35",x"f6",x"34",x"06",x"bd",x"f5",x"17",x"1f",
    x"89",x"84",x"30",x"a7",x"61",x"c4",x"0f",x"c1",x"04",x"24",x"02",x"cb",
    x"04",x"c1",x"0c",x"23",x"02",x"c0",x"04",x"eb",x"61",x"e7",x"61",x"35",
    x"86",x"34",x"06",x"86",x"7f",x"97",x"04",x"1f",x"20",x"bd",x"f2",x"c3",
    x"bd",x"f3",x"54",x"35",x"86",x"34",x"06",x"86",x"7f",x"97",x"04",x"a6",
    x"a4",x"e6",x"22",x"bd",x"f2",x"c3",x"bd",x"f3",x"54",x"35",x"86",x"34",
    x"16",x"1f",x"20",x"bd",x"f2",x"fc",x"e6",x"61",x"bd",x"f4",x"0e",x"35",
    x"96",x"34",x"16",x"1f",x"21",x"bd",x"f2",x"f2",x"e6",x"61",x"ae",x"62",
    x"bd",x"f4",x"0e",x"35",x"96",x"34",x"56",x"86",x"7f",x"97",x"04",x"bd",
    x"f3",x"73",x"35",x"d6",x"34",x"56",x"1f",x"20",x"bd",x"f2",x"fc",x"bd",
    x"f4",x"95",x"35",x"b6",x"bd",x"f2",x"a9",x"cc",x"fc",x"38",x"fd",x"c8",
    x"2a",x"b6",x"c8",x"9b",x"10",x"8e",x"ed",x"a3",x"10",x"ae",x"a6",x"ce",
    x"ed",x"9f",x"ee",x"c6",x"8d",x"da",x"39",x"bd",x"f2",x"a9",x"cc",x"fc",
    x"38",x"fd",x"c8",x"2a",x"10",x"8e",x"7f",x"a0",x"ce",x"c8",x"a8",x"8d",
    x"c7",x"b6",x"c8",x"79",x"27",x"09",x"10",x"8e",x"7f",x"10",x"ce",x"c8",
    x"af",x"8d",x"b9",x"39",x"bd",x"f1",x"92",x"34",x"08",x"bd",x"f2",x"e6",
    x"bd",x"ea",x"b4",x"b6",x"c8",x"80",x"bd",x"f1",x"b4",x"fc",x"c8",x"81",
    x"fd",x"c8",x"1f",x"fd",x"c8",x"21",x"bd",x"f1",x"f8",x"86",x"c8",x"1f",
    x"8b",x"96",x"9c",x"27",x"08",x"0a",x"9c",x"26",x"04",x"ad",x"9f",x"c8",
    x"9d",x"96",x"9f",x"27",x"08",x"0a",x"9f",x"26",x"04",x"ad",x"9f",x"c8",
    x"a0",x"96",x"a2",x"27",x"08",x"0a",x"a2",x"26",x"04",x"ad",x"9f",x"c8",
    x"a3",x"96",x"a5",x"27",x"08",x"0a",x"a5",x"26",x"04",x"ad",x"9f",x"c8",
    x"a6",x"35",x"88",x"96",x"ea",x"27",x"12",x"10",x"8e",x"c9",x"0b",x"86",
    x"04",x"97",x"8f",x"6d",x"a4",x"26",x"07",x"31",x"2a",x"0a",x"8f",x"26",
    x"f6",x"39",x"96",x"e7",x"27",x"35",x"34",x"20",x"a6",x"25",x"e6",x"27",
    x"1f",x"01",x"cc",x"06",x"16",x"10",x"9e",x"dc",x"bd",x"f8",x"ff",x"35",
    x"20",x"24",x"20",x"6f",x"a4",x"0f",x"e7",x"0f",x"a2",x"8e",x"ed",x"9f",
    x"96",x"9b",x"ae",x"86",x"cc",x"10",x"00",x"bd",x"f8",x"7c",x"86",x"30",
    x"c6",x"70",x"9e",x"dc",x"bd",x"e7",x"84",x"0a",x"ea",x"20",x"c6",x"ce",
    x"c9",x"33",x"86",x"1c",x"97",x"90",x"a6",x"c4",x"84",x"3f",x"26",x"09",
    x"33",x"c8",x"12",x"0a",x"90",x"26",x"f3",x"20",x"aa",x"34",x"20",x"a6",
    x"25",x"e6",x"27",x"1f",x"01",x"a6",x"44",x"e6",x"46",x"1f",x"02",x"ec",
    x"4c",x"bd",x"f8",x"ff",x"35",x"20",x"24",x"e0",x"a6",x"41",x"84",x"02",
    x"27",x"5a",x"8e",x"ed",x"9f",x"96",x"9b",x"ae",x"86",x"ec",x"4e",x"bd",
    x"f8",x"7c",x"0c",x"f5",x"a6",x"44",x"e6",x"46",x"1f",x"01",x"a6",x"42",
    x"c6",x"20",x"bd",x"e7",x"84",x"cc",x"01",x"10",x"ed",x"4e",x"96",x"c8",
    x"a0",x"44",x"d6",x"ca",x"e0",x"46",x"bd",x"f5",x"93",x"80",x"10",x"1f",
    x"89",x"34",x"20",x"86",x"3f",x"bd",x"e7",x"b5",x"10",x"af",x"48",x"af",
    x"4a",x"35",x"20",x"6f",x"a4",x"cc",x"04",x"04",x"ed",x"4c",x"a6",x"41",
    x"e6",x"43",x"5a",x"27",x"06",x"bd",x"e9",x"a1",x"bd",x"e9",x"a1",x"86",
    x"04",x"a7",x"41",x"0a",x"ea",x"7e",x"eb",x"53",x"86",x"01",x"a7",x"c4",
    x"6f",x"a4",x"8e",x"ed",x"9f",x"96",x"9b",x"ae",x"86",x"ec",x"4e",x"bd",
    x"f8",x"7c",x"a6",x"44",x"e6",x"46",x"1f",x"01",x"a6",x"42",x"c6",x"40",
    x"bd",x"e7",x"84",x"0a",x"eb",x"0a",x"ea",x"7e",x"eb",x"53",x"96",x"bd",
    x"26",x"19",x"96",x"ee",x"26",x"15",x"10",x"8e",x"c9",x"33",x"86",x"1c",
    x"97",x"8f",x"a6",x"a4",x"84",x"3f",x"26",x"08",x"31",x"a8",x"12",x"0a",
    x"8f",x"26",x"f3",x"39",x"34",x"20",x"96",x"c8",x"d6",x"ca",x"1f",x"01",
    x"a6",x"24",x"e6",x"26",x"10",x"ae",x"2c",x"1e",x"20",x"bd",x"f8",x"ff",
    x"35",x"20",x"24",x"e0",x"6f",x"a4",x"0f",x"ed",x"96",x"c8",x"d6",x"ca",
    x"1f",x"01",x"a6",x"22",x"8a",x"80",x"c6",x"30",x"bd",x"e7",x"84",x"0c",
    x"f3",x"0a",x"eb",x"20",x"ce",x"96",x"bd",x"26",x"19",x"96",x"ee",x"26",
    x"15",x"96",x"e7",x"27",x"11",x"96",x"c8",x"d6",x"ca",x"1f",x"01",x"cc",
    x"06",x"16",x"10",x"9e",x"dc",x"bd",x"f8",x"ff",x"25",x"01",x"39",x"0f",
    x"e7",x"0f",x"a2",x"96",x"c8",x"d6",x"ca",x"1f",x"01",x"86",x"08",x"8a",
    x"80",x"c6",x"30",x"bd",x"e7",x"84",x"0c",x"f3",x"39",x"b6",x"c8",x"f2",
    x"27",x"08",x"7f",x"c8",x"f2",x"ce",x"ed",x"37",x"20",x"31",x"b6",x"c8",
    x"f3",x"27",x"08",x"7f",x"c8",x"f3",x"ce",x"ed",x"4d",x"20",x"24",x"b6",
    x"c8",x"b6",x"27",x"08",x"7f",x"c8",x"b6",x"ce",x"ed",x"42",x"20",x"17",
    x"b6",x"c8",x"f4",x"27",x"0b",x"7f",x"c8",x"f4",x"7f",x"c8",x"f6",x"ce",
    x"ed",x"5a",x"20",x"07",x"b6",x"c8",x"f6",x"26",x"f0",x"20",x"03",x"bd",
    x"f2",x"7d",x"f6",x"c8",x"00",x"cb",x"10",x"c1",x"a0",x"24",x"07",x"86",
    x"00",x"bd",x"f2",x"56",x"20",x"06",x"cc",x"08",x"00",x"bd",x"f2",x"56",
    x"f6",x"c8",x"02",x"cb",x"20",x"c1",x"f0",x"24",x"07",x"86",x"02",x"bd",
    x"f2",x"56",x"20",x"06",x"cc",x"09",x"00",x"bd",x"f2",x"56",x"39",x"00",
    x"10",x"01",x"00",x"06",x"1f",x"07",x"06",x"08",x"0f",x"ff",x"02",x"39",
    x"03",x"00",x"06",x"1f",x"07",x"05",x"09",x"0f",x"ff",x"06",x"1f",x"07",
    x"07",x"0a",x"10",x"0b",x"00",x"0c",x"38",x"0d",x"00",x"ff",x"00",x"00",
    x"01",x"00",x"02",x"30",x"03",x"00",x"04",x"00",x"05",x"00",x"06",x"1f",
    x"07",x"3d",x"08",x"00",x"09",x"0f",x"0a",x"00",x"0b",x"00",x"0c",x"00",
    x"0d",x"00",x"ff",x"ed",x"8f",x"fe",x"b6",x"00",x"19",x"01",x"19",x"00",
    x"19",x"01",x"32",x"00",x"19",x"01",x"19",x"00",x"19",x"06",x"19",x"05",
    x"19",x"00",x"80",x"ff",x"ee",x"dd",x"cc",x"bb",x"aa",x"99",x"88",x"77",
    x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"c8",x"a8",x"c8",x"af",x"7f",
    x"a0",x"7f",x"10",x"c8",x"f9",x"c9",x"00",x"00",x"00",x"00",x"00",x"02",
    x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"02",
    x"01",x"00",x"00",x"02",x"03",x"00",x"00",x"01",x"03",x"00",x"00",x"02",
    x"02",x"00",x"00",x"01",x"01",x"00",x"00",x"03",x"03",x"00",x"00",x"02",
    x"02",x"02",x"00",x"01",x"01",x"01",x"00",x"03",x"03",x"03",x"00",x"80",
    x"c8",x"40",x"3f",x"00",x"20",x"80",x"10",x"1f",x"3f",x"3f",x"00",x"bf",
    x"bf",x"bf",x"c0",x"20",x"48",x"08",x"f8",x"30",x"a8",x"10",x"d0",x"a0",
    x"bf",x"bf",x"00",x"3f",x"3f",x"48",x"20",x"80",x"00",x"b0",x"48",x"38",
    x"fb",x"38",x"80",x"28",x"30",x"48",x"80",x"80",x"45",x"f0",x"28",x"7f",
    x"3f",x"bf",x"a5",x"00",x"d0",x"60",x"20",x"28",x"b8",x"40",x"15",x"80",
    x"40",x"f8",x"40",x"18",x"fa",x"38",x"e0",x"c8",x"4d",x"49",x"4e",x"45",
    x"20",x"46",x"49",x"45",x"4c",x"44",x"80",x"fa",x"38",x"e0",x"d8",x"47",
    x"41",x"4d",x"45",x"20",x"4f",x"56",x"45",x"52",x"80",x"00",x"10",x"00",
    x"ff",x"20",x"a0",x"ff",x"c0",x"40",x"ff",x"90",x"20",x"ff",x"70",x"20",
    x"ff",x"50",x"50",x"ff",x"d0",x"90",x"01",x"00",x"20",x"00",x"ff",x"30",
    x"b0",x"ff",x"b0",x"30",x"ff",x"b0",x"d0",x"ff",x"30",x"50",x"ff",x"d0",
    x"50",x"ff",x"50",x"d0",x"ff",x"50",x"30",x"ff",x"d0",x"b0",x"01",x"ff",
    x"00",x"00",x"00",x"30",x"00",x"ff",x"10",x"c0",x"ff",x"c0",x"10",x"ff",
    x"c0",x"f0",x"ff",x"10",x"40",x"ff",x"f0",x"40",x"ff",x"40",x"f0",x"ff",
    x"40",x"10",x"ff",x"f0",x"c0",x"01",x"ff",x"00",x"00",x"00",x"f0",x"d0",
    x"ff",x"c0",x"40",x"ff",x"20",x"00",x"ff",x"40",x"40",x"ff",x"00",x"e0",
    x"ff",x"40",x"c0",x"ff",x"e0",x"00",x"ff",x"c0",x"c0",x"ff",x"00",x"20",
    x"01",x"00",x"3f",x"00",x"ff",x"80",x"00",x"00",x"3f",x"3f",x"ff",x"00",
    x"80",x"01",x"ff",x"7f",x"20",x"00",x"c0",x"10",x"ff",x"c0",x"d0",x"ff",
    x"20",x"7f",x"00",x"e0",x"c0",x"ff",x"00",x"c0",x"ff",x"e0",x"30",x"00",
    x"c0",x"00",x"ff",x"60",x"cd",x"ff",x"a0",x"00",x"00",x"20",x"d0",x"ff",
    x"3c",x"30",x"ff",x"00",x"82",x"00",x"30",x"30",x"ff",x"d0",x"50",x"ff",
    x"20",x"f0",x"01",x"00",x"3f",x"00",x"ff",x"c4",x"08",x"ff",x"d8",x"d8",
    x"ff",x"20",x"00",x"00",x"00",x"40",x"ff",x"e0",x"00",x"ff",x"28",x"d8",
    x"ff",x"3c",x"08",x"01",x"00",x"3f",x"00",x"ff",x"c4",x"08",x"01",x"00",
    x"04",x"08",x"ff",x"d8",x"d8",x"ff",x"20",x"00",x"01",x"00",x"3f",x"00",
    x"ff",x"c4",x"f8",x"01",x"00",x"04",x"f8",x"ff",x"d8",x"28",x"ff",x"20",
    x"00",x"01",x"00",x"20",x"00",x"ff",x"00",x"d8",x"ff",x"d0",x"a8",x"ff",
    x"f0",x"40",x"ff",x"08",x"18",x"ff",x"18",x"f0",x"ff",x"f0",x"b8",x"00",
    x"10",x"48",x"ff",x"08",x"00",x"ff",x"e8",x"10",x"ff",x"f8",x"00",x"00",
    x"08",x"00",x"ff",x"00",x"06",x"00",x"10",x"fa",x"ff",x"08",x"00",x"ff",
    x"00",x"f0",x"00",x"10",x"18",x"ff",x"f0",x"08",x"01",x"00",x"20",x"00",
    x"ff",x"00",x"28",x"ff",x"d0",x"58",x"ff",x"f0",x"c0",x"ff",x"08",x"e8",
    x"ff",x"18",x"10",x"ff",x"f0",x"48",x"00",x"10",x"b8",x"ff",x"08",x"00",
    x"ff",x"e8",x"f0",x"ff",x"f8",x"00",x"ff",x"08",x"00",x"ff",x"00",x"fa",
    x"00",x"10",x"06",x"ff",x"08",x"00",x"ff",x"00",x"10",x"00",x"10",x"e8",
    x"ff",x"f0",x"f8",x"01",x"ff",x"00",x"d8",x"ff",x"e8",x"08",x"ff",x"00",
    x"40",x"ff",x"18",x"08",x"ff",x"00",x"d8",x"00",x"08",x"e0",x"ff",x"10",
    x"00",x"ff",x"00",x"40",x"ff",x"f0",x"00",x"ff",x"00",x"c0",x"01",x"00",
    x"18",x"00",x"ff",x"00",x"20",x"ff",x"c8",x"70",x"ff",x"10",x"a0",x"ff",
    x"00",x"a0",x"ff",x"ec",x"a4",x"ff",x"39",x"6d",x"ff",x"00",x"20",x"01",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"10",x"ce",x"cb",x"ea",x"bd",x"f1",x"8b",x"cc",
    x"73",x"21",x"10",x"b3",x"cb",x"fe",x"27",x"5c",x"fd",x"cb",x"fe",x"7c",
    x"c8",x"3b",x"8e",x"cb",x"eb",x"bd",x"f8",x"4f",x"bd",x"f1",x"af",x"dc",
    x"25",x"10",x"83",x"01",x"01",x"26",x"02",x"d7",x"56",x"57",x"c4",x"03",
    x"8e",x"f0",x"fd",x"e6",x"85",x"d7",x"29",x"c6",x"02",x"d7",x"24",x"ce",
    x"fd",x"0d",x"bd",x"f6",x"87",x"bd",x"f1",x"92",x"bd",x"f2",x"89",x"bd",
    x"f2",x"a9",x"b6",x"c8",x"26",x"ce",x"f1",x"0c",x"85",x"20",x"27",x"02",
    x"33",x"4c",x"bd",x"f3",x"85",x"8e",x"f0",x"e9",x"bd",x"f3",x"08",x"86",
    x"03",x"bd",x"f4",x"34",x"7a",x"c8",x"24",x"26",x"f3",x"b6",x"c8",x"25",
    x"81",x"01",x"23",x"b0",x"bd",x"f1",x"af",x"86",x"cc",x"97",x"29",x"cc", 
    x"f1",x"01",x"dd",x"39",x"0f",x"25",x"0f",x"26",x"ce",x"00",x"00",x"8e",
    x"f1",x"01",x"c6",x"0b",x"a6",x"c0",x"a1",x"80",x"27",x"0d",x"c1",x"01",
    x"27",x"04",x"c1",x"05",x"23",x"05",x"ce",x"e0",x"00",x"20",x"07",x"5a",
    x"26",x"ea",x"d7",x"39",x"d7",x"3a",x"0c",x"56",x"df",x"37",x"ee",x"c4",
    x"bd",x"f1",x"af",x"cc",x"f8",x"48",x"dd",x"2a",x"bd",x"f6",x"87",x"bd",
    x"f1",x"92",x"bd",x"f2",x"89",x"bd",x"f2",x"a9",x"cc",x"c0",x"c0",x"fe",
    x"c8",x"39",x"bd",x"f3",x"7a",x"b6",x"c8",x"3b",x"26",x"0c",x"4a",x"ce",
    x"cb",x"eb",x"a7",x"46",x"cc",x"68",x"d0",x"bd",x"f3",x"7a",x"fe",x"c8",
    x"37",x"33",x"42",x"bd",x"f3",x"85",x"b6",x"c8",x"56",x"26",x"c5",x"be",
    x"c8",x"25",x"8c",x"00",x"7d",x"23",x"bd",x"6e",x"41",x"40",x"d6",x"00",
    x"56",x"81",x"00",x"00",x"a9",x"7e",x"00",x"39",x"dc",x"8e",x"00",x"00",
    x"4a",x"72",x"00",x"00",x"b6",x"e0",x"38",x"0e",x"03",x"67",x"20",x"47",
    x"43",x"45",x"20",x"31",x"39",x"38",x"32",x"80",x"f1",x"60",x"27",x"cf",
    x"56",x"45",x"43",x"54",x"52",x"45",x"58",x"80",x"f3",x"60",x"26",x"cf",
    x"56",x"45",x"43",x"54",x"52",x"45",x"58",x"80",x"fc",x"60",x"df",x"e9",
    x"47",x"43",x"45",x"80",x"fc",x"38",x"cc",x"d1",x"45",x"4e",x"54",x"45",
    x"52",x"54",x"41",x"49",x"4e",x"49",x"4e",x"47",x"80",x"fc",x"38",x"bc",
    x"dc",x"4e",x"45",x"57",x"20",x"49",x"44",x"45",x"41",x"53",x"80",x"00",
    x"8d",x"5c",x"cc",x"9f",x"ff",x"dd",x"02",x"cc",x"01",x"00",x"dd",x"00",
    x"cc",x"98",x"7f",x"97",x"0b",x"d7",x"04",x"bd",x"f3",x"54",x"20",x"3e",
    x"8d",x"49",x"c6",x"7a",x"8e",x"c8",x"00",x"bd",x"f5",x"3f",x"cc",x"c8",
    x"7d",x"dd",x"7b",x"0c",x"7d",x"27",x"fc",x"86",x"05",x"97",x"28",x"cc",
    x"30",x"75",x"dd",x"3d",x"cc",x"01",x"03",x"dd",x"1f",x"cc",x"05",x"07",
    x"dd",x"21",x"39",x"8d",x"d7",x"8d",x"bd",x"7e",x"f2",x"72",x"be",x"c8",
    x"25",x"30",x"01",x"bf",x"c8",x"25",x"8d",x"0e",x"86",x"20",x"95",x"0d",
    x"27",x"fc",x"fc",x"c8",x"3d",x"dd",x"08",x"7e",x"f2",x"e6",x"86",x"d0",
    x"1f",x"8b",x"39",x"86",x"c8",x"1f",x"8b",x"39",x"b4",x"c8",x"0f",x"b7",
    x"c8",x"0f",x"8e",x"c8",x"12",x"a6",x"1d",x"a7",x"1e",x"86",x"0e",x"97",
    x"01",x"cc",x"19",x"01",x"97",x"00",x"12",x"d7",x"00",x"0f",x"03",x"cc",
    x"09",x"01",x"97",x"00",x"12",x"96",x"01",x"43",x"a7",x"1d",x"d7",x"00",
    x"c6",x"ff",x"d7",x"03",x"43",x"aa",x"1e",x"43",x"a7",x"1f",x"34",x"02",
    x"c6",x"01",x"1f",x"98",x"a4",x"e4",x"a7",x"80",x"58",x"26",x"f7",x"35",
    x"82",x"7a",x"c8",x"23",x"8e",x"c8",x"1f",x"a6",x"80",x"26",x"0c",x"8c",
    x"c8",x"23",x"26",x"f7",x"6f",x"84",x"86",x"01",x"97",x"00",x"39",x"97",
    x"00",x"0f",x"01",x"0a",x"00",x"c6",x"60",x"5c",x"2a",x"fd",x"b6",x"c8",
    x"23",x"2b",x"25",x"86",x"20",x"0c",x"00",x"95",x"00",x"27",x"0a",x"c6",
    x"40",x"d7",x"01",x"95",x"00",x"26",x"0b",x"20",x"08",x"c6",x"c0",x"d7",
    x"01",x"95",x"00",x"27",x"01",x"5f",x"e7",x"1b",x"20",x"c5",x"1f",x"98",
    x"9a",x"01",x"97",x"01",x"86",x"20",x"95",x"00",x"26",x"06",x"1f",x"98",
    x"98",x"01",x"97",x"01",x"54",x"f1",x"c8",x"1a",x"26",x"e8",x"d6",x"01",
    x"20",x"e0",x"8e",x"c8",x"00",x"e7",x"86",x"97",x"01",x"86",x"19",x"97",
    x"00",x"86",x"01",x"97",x"00",x"96",x"01",x"d7",x"01",x"c6",x"11",x"d7",
    x"00",x"c6",x"01",x"d7",x"00",x"39",x"cc",x"0e",x"00",x"8d",x"df",x"4a",
    x"2a",x"fb",x"7e",x"f5",x"33",x"8e",x"c8",x"00",x"20",x"02",x"8d",x"d5",
    x"ec",x"c1",x"2a",x"fa",x"39",x"8e",x"c8",x"00",x"ce",x"c8",x"3f",x"86",
    x"0d",x"e6",x"c0",x"e1",x"86",x"27",x"02",x"8d",x"c0",x"4a",x"2a",x"f5",
    x"39",x"86",x"1f",x"20",x"0a",x"86",x"3f",x"20",x"06",x"86",x"5f",x"20",
    x"02",x"86",x"7f",x"97",x"01",x"b7",x"c8",x"27",x"cc",x"05",x"04",x"97",
    x"00",x"d7",x"00",x"d7",x"00",x"c6",x"01",x"d7",x"00",x"39",x"f7",x"c8",
    x"28",x"ec",x"81",x"8d",x"4d",x"86",x"ff",x"97",x"0a",x"f6",x"c8",x"28",
    x"5a",x"26",x"fd",x"0f",x"0a",x"39",x"7a",x"c8",x"23",x"8d",x"ea",x"b6",
    x"c8",x"23",x"26",x"f6",x"20",x"76",x"a6",x"80",x"2e",x"72",x"8d",x"dd",
    x"20",x"f8",x"8e",x"f9",x"f0",x"8d",x"1d",x"bd",x"f3",x"6b",x"8d",x"20",
    x"20",x"62",x"c6",x"7f",x"d7",x"04",x"a6",x"84",x"e6",x"02",x"20",x"16",
    x"97",x"01",x"34",x"06",x"86",x"7f",x"97",x"04",x"0f",x"00",x"20",x"10",
    x"c6",x"ff",x"20",x"02",x"c6",x"7f",x"d7",x"04",x"ec",x"81",x"97",x"01",
    x"0f",x"00",x"34",x"06",x"86",x"ce",x"97",x"0c",x"0f",x"0a",x"0c",x"00",
    x"d7",x"01",x"0f",x"05",x"35",x"06",x"bd",x"f5",x"84",x"e7",x"7f",x"aa",
    x"7f",x"c6",x"40",x"81",x"40",x"23",x"12",x"81",x"64",x"23",x"04",x"86",
    x"08",x"20",x"02",x"86",x"04",x"d5",x"0d",x"27",x"fc",x"4a",x"26",x"fd",
    x"39",x"d5",x"0d",x"27",x"fc",x"39",x"bd",x"f1",x"aa",x"20",x"05",x"b6",
    x"c8",x"24",x"27",x"16",x"cc",x"00",x"cc",x"d7",x"0c",x"97",x"0a",x"cc",
    x"03",x"02",x"0f",x"01",x"97",x"00",x"d7",x"00",x"d7",x"00",x"c6",x"01",
    x"d7",x"00",x"39",x"cc",x"00",x"cc",x"d7",x"0c",x"97",x"0a",x"39",x"ec",
    x"c1",x"fd",x"c8",x"2a",x"ec",x"c1",x"bd",x"f2",x"fc",x"bd",x"f5",x"75",
    x"7e",x"f4",x"95",x"8d",x"ee",x"a6",x"c4",x"26",x"fa",x"39",x"8d",x"ec",
    x"a6",x"c4",x"26",x"fa",x"39",x"ae",x"84",x"34",x"04",x"c6",x"80",x"33",
    x"78",x"36",x"06",x"35",x"02",x"81",x"09",x"23",x"02",x"86",x"3c",x"8b",
    x"30",x"c6",x"2d",x"36",x"06",x"36",x"10",x"20",x"cb",x"a6",x"80",x"20",
    x"08",x"d7",x"04",x"20",x"07",x"ec",x"81",x"d7",x"04",x"b7",x"c8",x"23",
    x"ec",x"84",x"97",x"01",x"0f",x"00",x"30",x"02",x"12",x"0c",x"00",x"d7",
    x"01",x"cc",x"00",x"00",x"20",x"1f",x"a6",x"80",x"20",x"08",x"d7",x"04",
    x"20",x"07",x"ec",x"81",x"d7",x"04",x"b7",x"c8",x"23",x"ec",x"84",x"97",
    x"01",x"0f",x"00",x"30",x"02",x"12",x"0c",x"00",x"d7",x"01",x"cc",x"ff",
    x"00",x"97",x"0a",x"d7",x"05",x"cc",x"00",x"40",x"d5",x"0d",x"27",x"fc",
    x"12",x"97",x"0a",x"b6",x"c8",x"23",x"4a",x"2a",x"d9",x"7e",x"f3",x"4f",
    x"c6",x"ff",x"20",x"06",x"c6",x"7f",x"20",x"02",x"e6",x"80",x"d7",x"04",
    x"ec",x"01",x"97",x"01",x"0f",x"00",x"a6",x"84",x"30",x"03",x"0c",x"00",
    x"d7",x"01",x"97",x"0a",x"0f",x"05",x"cc",x"00",x"40",x"d5",x"0d",x"27",
    x"fc",x"12",x"97",x"0a",x"a6",x"84",x"2f",x"e0",x"7e",x"f3",x"4f",x"4a",
    x"b7",x"c8",x"23",x"ec",x"84",x"97",x"01",x"0f",x"00",x"30",x"02",x"0c",
    x"00",x"d7",x"01",x"b6",x"c8",x"29",x"c6",x"40",x"97",x"0a",x"0f",x"05",
    x"f5",x"d0",x"0d",x"27",x"0b",x"0f",x"0a",x"b6",x"c8",x"23",x"26",x"db",
    x"39",x"b6",x"c8",x"29",x"97",x"0a",x"12",x"d5",x"0d",x"27",x"f6",x"b6",
    x"c8",x"23",x"0f",x"0a",x"4d",x"26",x"c8",x"7e",x"f3",x"4f",x"b6",x"c8",
    x"24",x"34",x"02",x"7f",x"c8",x"24",x"a6",x"80",x"2a",x"04",x"8d",x"bb",
    x"20",x"f8",x"26",x"05",x"bd",x"f3",x"bc",x"20",x"f1",x"4a",x"27",x"05",
    x"bd",x"f3",x"dd",x"20",x"e9",x"35",x"02",x"b7",x"c8",x"24",x"7e",x"f3",
    x"4f",x"ff",x"c8",x"2c",x"8e",x"f9",x"d4",x"cc",x"18",x"83",x"0f",x"01",
    x"97",x"0b",x"8e",x"f9",x"d4",x"d7",x"00",x"0a",x"00",x"cc",x"80",x"81",
    x"12",x"0c",x"00",x"d7",x"00",x"97",x"00",x"7d",x"c8",x"00",x"0c",x"00",
    x"b6",x"c8",x"2b",x"97",x"01",x"cc",x"01",x"00",x"fe",x"c8",x"2c",x"97",
    x"00",x"20",x"04",x"a6",x"86",x"97",x"0a",x"a6",x"c0",x"2a",x"f8",x"86",
    x"81",x"97",x"00",x"00",x"01",x"86",x"01",x"97",x"00",x"8c",x"fb",x"b4",
    x"27",x"2c",x"30",x"88",x"50",x"1f",x"30",x"b3",x"c8",x"2c",x"c0",x"02",
    x"58",x"21",x"00",x"86",x"81",x"12",x"5a",x"26",x"fa",x"97",x"00",x"f6",
    x"c8",x"2a",x"d7",x"01",x"0a",x"00",x"cc",x"81",x"01",x"12",x"97",x"00",
    x"0f",x"01",x"d7",x"00",x"97",x"00",x"c6",x"03",x"20",x"9b",x"86",x"98",
    x"97",x"0b",x"7e",x"f3",x"54",x"34",x"14",x"c6",x"02",x"20",x"03",x"34",
    x"14",x"5f",x"be",x"c8",x"7b",x"a6",x"01",x"49",x"49",x"49",x"49",x"a8",
    x"02",x"46",x"69",x"84",x"69",x"01",x"69",x"02",x"5a",x"2a",x"ee",x"a6",
    x"84",x"35",x"94",x"c6",x"0d",x"8e",x"c8",x"3f",x"8d",x"05",x"86",x"3f",
    x"a7",x"06",x"39",x"4f",x"20",x"06",x"8e",x"c8",x"00",x"cc",x"00",x"ff",
    x"6f",x"8b",x"83",x"00",x"01",x"2a",x"f9",x"39",x"86",x"80",x"a7",x"85",
    x"5a",x"26",x"fb",x"a7",x"84",x"39",x"c6",x"02",x"20",x"02",x"c6",x"05",
    x"8e",x"c8",x"2e",x"6d",x"85",x"27",x"02",x"6a",x"85",x"5a",x"2a",x"f7",
    x"39",x"c6",x"03",x"20",x"09",x"c6",x"02",x"20",x"05",x"c6",x"01",x"20",
    x"01",x"5f",x"5a",x"2a",x"fd",x"39",x"8e",x"f9",x"dc",x"a6",x"86",x"39",
    x"4d",x"2a",x"04",x"40",x"28",x"01",x"4a",x"5d",x"2a",x"04",x"50",x"28",
    x"01",x"5a",x"39",x"34",x"10",x"dd",x"34",x"59",x"c6",x"00",x"59",x"49",
    x"59",x"58",x"d7",x"36",x"dc",x"34",x"8d",x"e0",x"97",x"34",x"d1",x"34",
    x"23",x"08",x"0c",x"36",x"1e",x"89",x"20",x"02",x"44",x"54",x"81",x"09",
    x"22",x"fa",x"dd",x"34",x"d6",x"36",x"8e",x"fc",x"24",x"e6",x"85",x"8e",
    x"fc",x"2c",x"a6",x"86",x"9b",x"35",x"8b",x"0a",x"c5",x"01",x"26",x"04",
    x"eb",x"86",x"20",x"03",x"5a",x"e0",x"86",x"d7",x"36",x"96",x"36",x"35",
    x"90",x"8b",x"10",x"8e",x"fc",x"6d",x"5f",x"85",x"20",x"27",x"02",x"c6",
    x"80",x"84",x"1f",x"81",x"10",x"26",x"01",x"5c",x"a6",x"86",x"39",x"34",
    x"10",x"96",x"36",x"8d",x"e6",x"dd",x"37",x"96",x"36",x"8d",x"de",x"dd",
    x"39",x"35",x"90",x"c0",x"10",x"d7",x"36",x"97",x"3b",x"8d",x"e8",x"8d",
    x"54",x"40",x"34",x"02",x"8d",x"55",x"35",x"84",x"b7",x"c8",x"36",x"f7",
    x"c8",x"23",x"34",x"08",x"bd",x"f1",x"af",x"8d",x"d2",x"20",x"18",x"b7",
    x"c8",x"36",x"34",x"08",x"bd",x"f1",x"af",x"97",x"23",x"8d",x"c4",x"a6",
    x"80",x"a7",x"c0",x"2f",x"06",x"0f",x"23",x"35",x"88",x"0a",x"23",x"a6",
    x"80",x"8d",x"26",x"a7",x"c4",x"a6",x"84",x"8d",x"1a",x"ab",x"c4",x"a7",
    x"c0",x"a6",x"1f",x"8d",x"12",x"a7",x"c4",x"a6",x"80",x"8d",x"12",x"a0",
    x"c4",x"a7",x"c0",x"96",x"23",x"2b",x"d4",x"26",x"dc",x"35",x"88",x"97",
    x"3b",x"dc",x"37",x"20",x"04",x"97",x"3b",x"dc",x"39",x"d7",x"3c",x"c5",
    x"01",x"27",x"04",x"96",x"3b",x"20",x"0a",x"d6",x"3b",x"2a",x"03",x"03",
    x"3c",x"50",x"3d",x"89",x"00",x"d6",x"3c",x"2a",x"01",x"40",x"39",x"e6",
    x"c6",x"e7",x"86",x"4a",x"2a",x"f9",x"39",x"96",x"56",x"2b",x"28",x"27",
    x"f9",x"8e",x"fc",x"8d",x"9f",x"4d",x"86",x"80",x"97",x"56",x"ec",x"c1",
    x"dd",x"4f",x"ec",x"c1",x"dd",x"51",x"df",x"53",x"bd",x"f5",x"33",x"cc",
    x"1f",x"1f",x"dd",x"5f",x"cc",x"00",x"00",x"dd",x"63",x"dd",x"65",x"97",
    x"55",x"20",x"39",x"ce",x"c8",x"5e",x"c6",x"02",x"a6",x"c5",x"81",x"1f",
    x"27",x"02",x"6c",x"c5",x"5a",x"2a",x"f5",x"9e",x"51",x"ce",x"c8",x"58",
    x"86",x"07",x"6c",x"c4",x"a1",x"c4",x"2c",x"02",x"6f",x"c4",x"e6",x"c0",
    x"c4",x"07",x"e6",x"85",x"e7",x"c0",x"4c",x"81",x"09",x"23",x"eb",x"0a",
    x"57",x"26",x"6b",x"96",x"55",x"4a",x"2a",x"02",x"86",x"02",x"97",x"55",
    x"e6",x"9f",x"c8",x"53",x"ce",x"c8",x"5e",x"6f",x"c6",x"c5",x"40",x"27",
    x"19",x"8e",x"f9",x"e4",x"a6",x"86",x"94",x"45",x"97",x"45",x"96",x"55",
    x"8b",x"03",x"a6",x"86",x"9a",x"45",x"97",x"45",x"c4",x"1f",x"d7",x"46",
    x"20",x"23",x"8e",x"f9",x"ea",x"a6",x"86",x"94",x"45",x"97",x"45",x"96",
    x"55",x"8b",x"03",x"a6",x"86",x"9a",x"45",x"97",x"45",x"96",x"55",x"48",
    x"8b",x"03",x"33",x"c6",x"c4",x"3f",x"58",x"9e",x"4d",x"ec",x"85",x"ed",
    x"c4",x"9e",x"53",x"e6",x"80",x"9f",x"53",x"5d",x"2b",x"a5",x"e6",x"80",
    x"2a",x"06",x"bd",x"f5",x"33",x"0f",x"56",x"39",x"9f",x"53",x"c4",x"3f",
    x"d7",x"57",x"10",x"9e",x"4f",x"ce",x"c8",x"5e",x"8e",x"c8",x"42",x"86",
    x"02",x"e6",x"c0",x"c5",x"01",x"27",x"07",x"54",x"e6",x"a5",x"c4",x"0f",
    x"20",x"07",x"54",x"e6",x"a5",x"54",x"54",x"54",x"54",x"e7",x"86",x"4a",
    x"2a",x"e7",x"ce",x"c8",x"67",x"8e",x"c8",x"47",x"ec",x"c3",x"6d",x"58",
    x"2a",x"0a",x"60",x"58",x"e0",x"58",x"82",x"00",x"60",x"58",x"20",x"04",
    x"eb",x"58",x"89",x"00",x"ed",x"81",x"8c",x"c8",x"4d",x"26",x"e5",x"39",
    x"20",x"c0",x"40",x"c0",x"50",x"4c",x"41",x"59",x"45",x"52",x"80",x"e0",
    x"c0",x"01",x"c0",x"20",x"47",x"41",x"4d",x"45",x"80",x"fd",x"c8",x"4f",
    x"4d",x"27",x"02",x"86",x"01",x"5d",x"27",x"02",x"c6",x"01",x"fd",x"c8",
    x"79",x"bd",x"f1",x"af",x"cc",x"f8",x"50",x"dd",x"2a",x"97",x"3c",x"20",
    x"67",x"bd",x"f1",x"92",x"4f",x"bd",x"f1",x"b4",x"bd",x"f5",x"5a",x"bd",
    x"f2",x"a9",x"b6",x"c8",x"79",x"10",x"8e",x"f7",x"94",x"8d",x"5a",x"b6",
    x"c8",x"7a",x"10",x"8e",x"f7",x"9f",x"8d",x"51",x"bd",x"f1",x"af",x"96",
    x"3c",x"27",x"06",x"96",x"0f",x"26",x"3d",x"0f",x"3c",x"96",x"2f",x"27",
    x"9e",x"96",x"2e",x"26",x"cc",x"96",x"15",x"26",x"96",x"96",x"12",x"27",
    x"0f",x"96",x"79",x"27",x"0b",x"4c",x"91",x"4f",x"23",x"02",x"86",x"01",
    x"97",x"79",x"20",x"1c",x"96",x"7a",x"27",x"b1",x"d6",x"13",x"27",x"09",
    x"4c",x"91",x"50",x"23",x"0d",x"86",x"01",x"20",x"09",x"d6",x"14",x"27",
    x"a0",x"4a",x"26",x"02",x"96",x"50",x"97",x"7a",x"86",x"f3",x"97",x"2f",
    x"43",x"97",x"2e",x"20",x"90",x"8e",x"c8",x"5e",x"34",x"02",x"8d",x"13",
    x"a6",x"e0",x"27",x"0e",x"8d",x"1c",x"1f",x"13",x"ec",x"a1",x"bd",x"f3",
    x"7a",x"1f",x"23",x"bd",x"f3",x"78",x"39",x"cc",x"20",x"20",x"ed",x"84",
    x"ed",x"02",x"a7",x"04",x"cc",x"30",x"80",x"ed",x"05",x"39",x"ce",x"00",
    x"00",x"81",x"63",x"23",x"08",x"80",x"64",x"33",x"c9",x"01",x"00",x"20",
    x"f4",x"81",x"09",x"23",x"07",x"80",x"0a",x"33",x"c8",x"10",x"20",x"f5",
    x"33",x"c6",x"1f",x"30",x"34",x"02",x"34",x"04",x"c6",x"05",x"4f",x"c1",
    x"01",x"23",x"10",x"c5",x"01",x"27",x"04",x"a6",x"e4",x"20",x"06",x"a6",
    x"e0",x"44",x"44",x"44",x"44",x"84",x"0f",x"bb",x"c8",x"23",x"7f",x"c8",
    x"23",x"ab",x"85",x"81",x"2f",x"2e",x"02",x"8b",x"10",x"81",x"39",x"23",
    x"05",x"80",x"0a",x"7c",x"c8",x"23",x"a7",x"85",x"5a",x"2a",x"cf",x"7f",
    x"c8",x"23",x"5f",x"a6",x"85",x"81",x"30",x"26",x"09",x"86",x"20",x"a7",
    x"85",x"5c",x"c1",x"05",x"2d",x"f1",x"39",x"34",x"50",x"4f",x"e6",x"80",
    x"2b",x"08",x"e1",x"c0",x"27",x"f8",x"22",x"01",x"4c",x"4c",x"35",x"d0",
    x"8d",x"ed",x"81",x"01",x"26",x"06",x"a6",x"80",x"a7",x"c0",x"2a",x"fa",
    x"39",x"34",x"20",x"34",x"36",x"ec",x"64",x"ab",x"c4",x"eb",x"41",x"ed",
    x"64",x"20",x"10",x"34",x"20",x"34",x"36",x"1f",x"30",x"ab",x"64",x"eb",
    x"65",x"20",x"f0",x"34",x"20",x"34",x"36",x"1f",x"41",x"5f",x"3a",x"a6",
    x"04",x"ab",x"84",x"28",x"02",x"86",x"7f",x"a1",x"02",x"2d",x"15",x"a6",
    x"04",x"a0",x"84",x"28",x"02",x"86",x"80",x"a1",x"02",x"2e",x"09",x"5c",
    x"c1",x"02",x"25",x"e2",x"1a",x"01",x"20",x"02",x"1c",x"fe",x"35",x"36",
    x"35",x"a0",x"96",x"67",x"2a",x"29",x"84",x"7f",x"97",x"67",x"8e",x"c8",
    x"58",x"86",x"04",x"bd",x"f6",x"83",x"54",x"54",x"54",x"da",x"58",x"c4",
    x"07",x"d7",x"54",x"d6",x"58",x"c4",x"38",x"d7",x"53",x"d6",x"58",x"c4",
    x"07",x"d7",x"5d",x"c6",x"02",x"d7",x"5c",x"86",x"7f",x"20",x"0d",x"96",
    x"77",x"27",x"6a",x"90",x"5b",x"2a",x"05",x"5f",x"d7",x"77",x"20",x"62",
    x"97",x"77",x"44",x"44",x"d6",x"53",x"27",x"0d",x"97",x"46",x"d6",x"59",
    x"2b",x"05",x"27",x"05",x"1f",x"89",x"53",x"d7",x"46",x"44",x"81",x"07",
    x"23",x"05",x"81",x"0f",x"27",x"01",x"4c",x"d6",x"5a",x"2b",x"06",x"27",
    x"02",x"88",x"0f",x"1f",x"89",x"8d",x"37",x"d6",x"5d",x"27",x"2b",x"96",
    x"5c",x"4a",x"2a",x"02",x"86",x"02",x"97",x"5c",x"bd",x"f5",x"7e",x"95",
    x"5d",x"27",x"f0",x"d6",x"5c",x"58",x"50",x"8e",x"c8",x"4b",x"30",x"85",
    x"bd",x"f5",x"17",x"84",x"0f",x"81",x"05",x"22",x"03",x"48",x"8b",x"05",
    x"a7",x"84",x"96",x"7e",x"a7",x"01",x"96",x"58",x"43",x"94",x"45",x"97",
    x"45",x"39",x"96",x"54",x"8e",x"c8",x"45",x"4d",x"27",x"09",x"30",x"1f",
    x"44",x"24",x"f8",x"e7",x"84",x"20",x"f4",x"39",x"01",x"02",x"04",x"08",
    x"10",x"20",x"40",x"80",x"f7",x"ef",x"df",x"01",x"02",x"04",x"fe",x"fd",
    x"fb",x"08",x"10",x"20",x"7f",x"7f",x"80",x"80",x"00",x"20",x"50",x"50",
    x"20",x"c8",x"20",x"10",x"10",x"40",x"20",x"00",x"00",x"00",x"00",x"08",
    x"30",x"20",x"70",x"70",x"10",x"f8",x"30",x"f8",x"70",x"70",x"00",x"60",
    x"00",x"00",x"00",x"70",x"70",x"20",x"f0",x"70",x"f0",x"f8",x"f8",x"78",
    x"88",x"70",x"08",x"88",x"80",x"88",x"88",x"f8",x"f0",x"70",x"f0",x"70",
    x"f8",x"88",x"88",x"88",x"88",x"88",x"f8",x"70",x"80",x"70",x"20",x"00",
    x"00",x"20",x"08",x"20",x"00",x"00",x"00",x"38",x"10",x"20",x"44",x"44",
    x"00",x"fe",x"ff",x"fe",x"00",x"70",x"50",x"50",x"78",x"c8",x"50",x"20",
    x"20",x"20",x"a8",x"20",x"00",x"00",x"00",x"08",x"48",x"60",x"88",x"88",
    x"30",x"80",x"40",x"08",x"88",x"88",x"60",x"60",x"10",x"00",x"40",x"88",
    x"88",x"50",x"48",x"88",x"48",x"80",x"80",x"80",x"88",x"20",x"08",x"90",
    x"80",x"d8",x"c8",x"88",x"88",x"88",x"88",x"88",x"a8",x"88",x"88",x"88",
    x"88",x"88",x"08",x"40",x"80",x"08",x"50",x"00",x"00",x"70",x"0c",x"20",
    x"70",x"70",x"00",x"44",x"10",x"70",x"00",x"00",x"6c",x"82",x"ff",x"fe",
    x"00",x"70",x"50",x"f8",x"a0",x"10",x"50",x"40",x"40",x"10",x"70",x"20",
    x"00",x"00",x"00",x"10",x"48",x"20",x"08",x"08",x"50",x"f0",x"80",x"10",
    x"88",x"88",x"60",x"00",x"20",x"78",x"20",x"08",x"a8",x"88",x"48",x"80",
    x"48",x"80",x"80",x"80",x"88",x"20",x"08",x"a0",x"80",x"a8",x"a8",x"88",
    x"88",x"88",x"88",x"40",x"20",x"88",x"88",x"88",x"50",x"50",x"10",x"40",
    x"40",x"08",x"88",x"00",x"70",x"a8",x"0a",x"20",x"88",x"f8",x"60",x"ba",
    x"38",x"20",x"00",x"00",x"92",x"82",x"ff",x"fe",x"00",x"20",x"00",x"50",
    x"70",x"20",x"60",x"00",x"40",x"10",x"a8",x"f8",x"00",x"70",x"00",x"20",
    x"48",x"20",x"70",x"30",x"90",x"08",x"f0",x"20",x"70",x"78",x"00",x"60",
    x"40",x"00",x"10",x"10",x"b8",x"88",x"70",x"80",x"48",x"e0",x"e0",x"98",
    x"f8",x"20",x"08",x"c0",x"80",x"a8",x"98",x"88",x"f0",x"88",x"f0",x"20",
    x"20",x"88",x"50",x"a8",x"20",x"20",x"20",x"40",x"20",x"08",x"00",x"00",
    x"fe",x"20",x"08",x"20",x"88",x"f8",x"f0",x"a2",x"38",x"f8",x"82",x"38",
    x"92",x"82",x"ff",x"fe",x"00",x"00",x"00",x"f8",x"70",x"40",x"a8",x"00",
    x"40",x"10",x"a8",x"20",x"40",x"00",x"00",x"40",x"48",x"20",x"80",x"08",
    x"f8",x"08",x"88",x"40",x"88",x"08",x"60",x"60",x"20",x"78",x"20",x"20",
    x"b0",x"f8",x"48",x"80",x"48",x"80",x"80",x"88",x"88",x"20",x"08",x"a0",
    x"80",x"88",x"88",x"88",x"80",x"a8",x"a0",x"10",x"20",x"88",x"50",x"a8",
    x"50",x"20",x"40",x"40",x"10",x"08",x"00",x"00",x"fe",x"20",x"78",x"a8",
    x"88",x"f8",x"f0",x"ba",x"7c",x"20",x"44",x"44",x"6c",x"82",x"ff",x"fe",
    x"00",x"00",x"00",x"50",x"28",x"98",x"90",x"00",x"20",x"20",x"00",x"20",
    x"40",x"00",x"00",x"80",x"48",x"20",x"80",x"88",x"10",x"88",x"88",x"80",
    x"88",x"10",x"60",x"20",x"10",x"00",x"40",x"00",x"80",x"88",x"48",x"88",
    x"48",x"80",x"80",x"88",x"88",x"20",x"88",x"90",x"88",x"88",x"88",x"88",
    x"80",x"90",x"90",x"88",x"20",x"88",x"20",x"a8",x"88",x"20",x"80",x"40",
    x"08",x"08",x"00",x"00",x"48",x"20",x"f0",x"70",x"70",x"70",x"60",x"44",
    x"6c",x"50",x"38",x"82",x"00",x"82",x"ff",x"fe",x"00",x"20",x"00",x"50",
    x"f8",x"98",x"68",x"00",x"10",x"40",x"00",x"00",x"80",x"00",x"80",x"80",
    x"30",x"70",x"f8",x"70",x"10",x"70",x"70",x"80",x"70",x"60",x"00",x"40",
    x"00",x"00",x"00",x"20",x"78",x"88",x"f0",x"70",x"f0",x"f8",x"80",x"78",
    x"88",x"70",x"70",x"88",x"f8",x"88",x"88",x"f8",x"80",x"68",x"88",x"70",
    x"20",x"70",x"20",x"50",x"88",x"20",x"f8",x"70",x"08",x"70",x"00",x"f8",
    x"00",x"20",x"60",x"20",x"00",x"00",x"00",x"38",x"82",x"88",x"00",x"00",
    x"00",x"fe",x"ff",x"fe",x"00",x"11",x"41",x"30",x"21",x"10",x"20",x"31",
    x"00",x"01",x"03",x"06",x"0a",x"0f",x"15",x"1c",x"24",x"2d",x"08",x"10",
    x"08",x"10",x"0b",x"08",x"10",x"0d",x"0a",x"08",x"10",x"0e",x"0b",x"09",
    x"08",x"10",x"0e",x"0c",x"0a",x"09",x"08",x"10",x"0e",x"0d",x"0b",x"0a",
    x"09",x"08",x"10",x"0f",x"0d",x"0c",x"0b",x"0a",x"09",x"08",x"10",x"0f",
    x"0e",x"0c",x"0b",x"0a",x"09",x"09",x"08",x"10",x"0f",x"0e",x"0d",x"0c",
    x"0b",x"0a",x"09",x"09",x"08",x"00",x"19",x"32",x"4a",x"62",x"79",x"8e",
    x"a2",x"b5",x"c6",x"d5",x"e2",x"ed",x"f5",x"fb",x"ff",x"ff",x"ff",x"fb",
    x"f5",x"ed",x"e2",x"d5",x"c6",x"b5",x"a2",x"8e",x"79",x"62",x"4a",x"32",
    x"19",x"03",x"bd",x"03",x"87",x"03",x"54",x"03",x"24",x"02",x"f7",x"02",
    x"cd",x"02",x"a4",x"02",x"7e",x"02",x"5b",x"02",x"39",x"02",x"19",x"01",
    x"fb",x"01",x"de",x"01",x"c3",x"01",x"aa",x"01",x"92",x"01",x"7c",x"01",
    x"66",x"01",x"52",x"01",x"3f",x"01",x"2d",x"01",x"1c",x"01",x"0c",x"00",
    x"fd",x"00",x"ef",x"00",x"e2",x"00",x"d5",x"00",x"c9",x"00",x"be",x"00",
    x"b3",x"00",x"a9",x"00",x"a0",x"00",x"97",x"00",x"8e",x"00",x"86",x"00",
    x"7f",x"00",x"78",x"00",x"71",x"00",x"6b",x"00",x"65",x"00",x"5f",x"00",
    x"5a",x"00",x"55",x"00",x"50",x"00",x"4b",x"00",x"47",x"00",x"43",x"00",
    x"3f",x"00",x"3c",x"00",x"38",x"00",x"35",x"00",x"32",x"00",x"2f",x"00",
    x"2d",x"00",x"2a",x"00",x"28",x"00",x"26",x"00",x"24",x"00",x"22",x"00",
    x"20",x"00",x"1e",x"00",x"1c",x"00",x"1b",x"00",x"00",x"fe",x"e8",x"fe",
    x"b6",x"93",x"1f",x"0c",x"93",x"1f",x"06",x"98",x"9f",x"24",x"3c",x"11",
    x"80",x"fd",x"69",x"fd",x"79",x"21",x"07",x"21",x"07",x"21",x"07",x"21",
    x"07",x"21",x"07",x"21",x"07",x"21",x"0e",x"99",x"9f",x"24",x"0e",x"95",
    x"9b",x"20",x"0e",x"21",x"07",x"21",x"07",x"21",x"07",x"21",x"07",x"21",
    x"07",x"21",x"07",x"9d",x"a3",x"28",x"0e",x"a0",x"a6",x"2b",x"0e",x"22",
    x"02",x"28",x"02",x"2d",x"02",x"28",x"02",x"22",x"02",x"28",x"02",x"2d",
    x"02",x"28",x"02",x"22",x"02",x"28",x"02",x"2d",x"02",x"28",x"02",x"2e",
    x"02",x"2d",x"28",x"21",x"80",x"ef",x"ff",x"fe",x"dc",x"ba",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",
    x"01",x"00",x"ff",x"fe",x"ff",x"fd",x"c3",x"fe",x"b6",x"51",x"24",x"50",
    x"06",x"50",x"06",x"50",x"0c",x"50",x"06",x"50",x"06",x"50",x"04",x"50",
    x"04",x"50",x"04",x"50",x"18",x"50",x"04",x"50",x"04",x"50",x"04",x"50",
    x"0c",x"50",x"0c",x"50",x"24",x"50",x"06",x"50",x"06",x"50",x"0c",x"50",
    x"06",x"50",x"06",x"50",x"04",x"50",x"04",x"50",x"04",x"50",x"18",x"50",
    x"04",x"50",x"04",x"50",x"04",x"50",x"0c",x"50",x"18",x"26",x"80",x"fd",
    x"ba",x"98",x"76",x"55",x"44",x"33",x"22",x"11",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"fe",x"28",x"fd",x"79",x"98",x"1c",x"10",x"3f",x"08",
    x"98",x"1c",x"04",x"98",x"1c",x"04",x"98",x"1c",x"10",x"3f",x"08",x"98",
    x"1c",x"04",x"98",x"1c",x"04",x"98",x"1c",x"08",x"93",x"18",x"08",x"98",
    x"1c",x"08",x"9c",x"1f",x"08",x"98",x"1c",x"08",x"93",x"18",x"08",x"98",
    x"1c",x"08",x"93",x"18",x"08",x"98",x"1c",x"08",x"9c",x"1f",x"08",x"98",
    x"1c",x"08",x"93",x"18",x"08",x"98",x"1c",x"08",x"93",x"18",x"08",x"98",
    x"1c",x"08",x"9c",x"1f",x"08",x"98",x"1c",x"08",x"93",x"18",x"08",x"9c",
    x"1f",x"30",x"1a",x"80",x"ff",x"fe",x"dc",x"ba",x"98",x"76",x"54",x"32",
    x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"66",x"fe",x"b6",
    x"0c",x"18",x"11",x"18",x"0c",x"18",x"11",x"18",x"0c",x"18",x"11",x"18",
    x"0c",x"12",x"0c",x"06",x"11",x"18",x"9d",x"21",x"18",x"9f",x"23",x"18",
    x"a1",x"24",x"18",x"a3",x"26",x"18",x"9f",x"a4",x"28",x"18",x"07",x"12",
    x"07",x"06",x"00",x"3c",x"18",x"80",x"de",x"ef",x"fe",x"dc",x"ba",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"b2",
    x"fe",x"b6",x"18",x"06",x"1a",x"06",x"1c",x"0c",x"18",x"0c",x"1a",x"24",
    x"23",x"18",x"17",x"06",x"18",x"06",x"1a",x"0c",x"17",x"0c",x"18",x"24",
    x"24",x"18",x"a4",x"28",x"0c",x"a3",x"26",x"0c",x"a1",x"24",x"0c",x"9f",
    x"23",x"0c",x"9d",x"21",x"18",x"9a",x"1f",x"18",x"17",x"06",x"18",x"06",
    x"1a",x"0c",x"17",x"0c",x"18",x"24",x"24",x"24",x"18",x"80",x"ff",x"ee",
    x"dd",x"cc",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"e8",x"fe",x"b6",x"96",x"9a",
    x"1d",x"1e",x"91",x"95",x"18",x"1e",x"94",x"98",x"1b",x"1e",x"8f",x"94",
    x"18",x"14",x"16",x"0a",x"8c",x"91",x"15",x"14",x"16",x"0a",x"91",x"95",
    x"18",x"32",x"18",x"80",x"ee",x"ff",x"ff",x"ee",x"ee",x"dd",x"cc",x"bb",
    x"aa",x"99",x"88",x"88",x"88",x"88",x"88",x"88",x"ff",x"16",x"fe",x"b6",
    x"1c",x"06",x"1f",x"06",x"1c",x"06",x"18",x"06",x"1a",x"06",x"18",x"06",
    x"15",x"06",x"13",x"06",x"18",x"06",x"13",x"06",x"17",x"06",x"18",x"1e",
    x"18",x"80",x"ff",x"ff",x"ee",x"ee",x"dd",x"dd",x"cc",x"cc",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"fe",x"28",x"fe",x"b6",x"16",x"0f",
    x"16",x"05",x"16",x"05",x"16",x"05",x"1a",x"0f",x"16",x"0f",x"1d",x"0f",
    x"1d",x"05",x"1d",x"05",x"1d",x"05",x"21",x"0f",x"1d",x"32",x"1d",x"80",
    x"fe",x"28",x"fe",x"b6",x"16",x"06",x"16",x"02",x"16",x"02",x"16",x"02",
    x"1a",x"06",x"16",x"06",x"1d",x"06",x"1d",x"02",x"1d",x"02",x"1d",x"02",
    x"21",x"06",x"1d",x"32",x"11",x"80",x"fe",x"28",x"fe",x"b6",x"1b",x"0f",
    x"16",x"05",x"16",x"05",x"16",x"05",x"17",x"30",x"16",x"05",x"16",x"05",
    x"16",x"05",x"17",x"30",x"16",x"80",x"fd",x"69",x"fe",x"b6",x"a0",x"23",
    x"12",x"a0",x"23",x"0c",x"9c",x"20",x"06",x"9e",x"21",x"12",x"9c",x"20",
    x"32",x"13",x"80",x"fd",x"c3",x"fe",x"b6",x"16",x"04",x"16",x"04",x"16",
    x"04",x"16",x"04",x"1a",x"08",x"1c",x"80",x"a6",x"a0",x"20",x"08",x"bd",
    x"f3",x"be",x"b6",x"c8",x"80",x"84",x"7f",x"b7",x"c8",x"80",x"7a",x"c8",
    x"80",x"a6",x"a4",x"47",x"84",x"f8",x"e6",x"a0",x"58",x"58",x"58",x"58",
    x"57",x"c4",x"f8",x"7d",x"c8",x"80",x"2b",x"df",x"bd",x"f3",x"df",x"b6",
    x"c8",x"80",x"85",x"0f",x"26",x"e0",x"85",x"20",x"27",x"cd",x"39",x"4b",
    x"41",x"52",x"52",x"53",x"4f",x"46",x"54",x"38",x"32",x"4c",x"44",x"4d",
    x"43",x"42",x"43",x"4a",x"54",x"38",x"32",x"4c",x"44",x"4d",x"43",x"42",
    x"43",x"4a",x"00",x"00",x"00",x"00",x"cb",x"f2",x"cb",x"f2",x"cb",x"f5",
    x"cb",x"f8",x"cb",x"fb",x"cb",x"fb",x"f0",x"00");

BEGIN
  PROCESS(clk) IS
  BEGIN
    IF rising_edge(clk) THEN
      dr<=rom(to_integer(ad AND x"1FFF"));
    END IF;
  END PROCESS;


  
    
END ARCHITECTURE rtl;

